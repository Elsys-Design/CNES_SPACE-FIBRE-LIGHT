----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module describe the Data_word_id_fsm function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_crc_check is
  port (
    RST_N              : in  std_logic;                                    --! global reset
    CLK                : in  std_logic;                                    --! Clock generated by GTY IP
    -- DWI interface
    DATA_DWI           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    NEW_WORD_DWI       : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    END_FRAME_DWI      : in  std_logic;
    SEQ_NUM_DWI        : in  std_logic_vector(7 downto 0);
    CRC_16B_DWI        : in  std_logic_vector(15 downto 0);                --! Flag EMPTY of the FIFO RX
    CRC_8B_DWI         : in  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
    TYPE_FRAME_DWI     : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);                 --! Flag EMPTY of the FIFO RX
    -- DWI interface
    NEW_WORD_DCCHECK   : out std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    DATA_DCCHECK       : out std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    END_FRAME_DCCHECK  : out std_logic;
    TYPE_FRAME_DCCHECK : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);                 --! Flag EMPTY of the FIFO RX
    SEQ_NUM_DCCHECK    : out std_logic_vector(7 downto 0);
    CRC_ERR            : out std_logic

  );
end data_crc_check;

architecture rtl of data_crc_check is

----------------------------- Declaration signals -----------------------------
type int_array     is array (0 to 3) of integer;
signal indices     : int_array := (0, 8, 16, 24);

type int_array_tier     is array (0 to 2) of integer;
signal indices_tier : int_array_tier := (0, 8, 16);

type int_array_dem is array (0 to 1) of integer;
signal indices_dem : int_array_dem := (0, 8);


signal crc_reg         : std_logic_vector(16-1 downto 0);   --! Data parallel from Lane Layer
signal crc_to_inv      : std_logic;                         --! Data parallel from Lane Layer
signal end_crc         : std_logic;                         --! Data parallel from Lane Layer
signal crc_err_16b     : std_logic;                         --! Data parallel from Lane Layer

signal crc_reg_8b      : std_logic_vector(8-1 downto 0);   --! Data parallel from Lane Layer
signal crc_to_inv_8b   : std_logic;                        --! Data parallel from Lane Layer
signal end_CRC_8B_DWI  : std_logic;                        --! Data parallel from Lane Layer
signal crc_err_8b      : std_logic;                        --! Data parallel from Lane Layer

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_CRC_16B_DWI
-- Description: Compute the CRC for a data frame 
---------------------------------------------------------
 p_CRC_16B_DWI: process(CLK, RST_N)
    variable crc_var : std_logic_vector(15 downto 0);
begin
    if RST_N = '0' then
        crc_reg        <= (others => '1'); -- Reset CRC to seed value
        crc_to_inv     <= '0';
        crc_err_16b    <= '0';
        end_crc        <= '0';
    elsif rising_edge(CLK) then
      crc_var := crc_reg;
      crc_err_16b    <= '0';
      if (TYPE_FRAME_DWI = C_DATA_FRM) then
        if end_crc = '1' then
          end_crc <= '0';
          if crc_reg /= CRC_16B_DWI then
            crc_err_16b <= '1';
          end if;
          crc_reg    <= (others => '1'); 

        elsif crc_to_inv = '1' then -- 
          crc_to_inv <= '0';
          end_crc    <= '1'; 
          for i in 0 to 15 loop
            crc_var(i) := crc_reg(15 - i); -- Bit-by-bit inversion
          end loop;
          crc_reg <= crc_var; 

        elsif END_FRAME_DWI = '1' and NEW_WORD_DWI = '1'then -- EDF detection
          crc_to_inv <= '1';
          for i in indices_dem'range loop -- calculates the crc 8 byte by byte
              crc_var := calculate_crc_16(DATA_DWI(7+ indices_dem(i) downto 0 + indices_dem(i)), crc_var);
          end loop;
          crc_reg <= crc_var; 

        elsif NEW_WORD_DWI = '1' then
          for i in indices'range loop -- calculates the crc 8 byte by byte
              crc_var := calculate_crc_16(DATA_DWI(7+ indices(i) downto 0 + indices(i)), crc_var);
          end loop;
          crc_reg <= crc_var; 
        end if;
      end if;
    end if;
end process p_CRC_16B_DWI;

---------------------------------------------------------
-- Process: p_CRC_8B_DWI
-- Description: Compute the CRC for broadcast frame, 
--              FCT, ACK, NACK and SIF
---------------------------------------------------------
p_CRC_8B_DWI: process(CLK, RST_N)
    variable crc_var : std_logic_vector(7 downto 0);
begin
    if RST_N = '0' then
        crc_reg_8b    <= (others => '0'); -- Reset CRC to seed value
        crc_to_inv_8b <= '0';
        crc_err_8b    <= '0';
        end_CRC_8B_DWI    <= '0';
    elsif rising_edge(CLK) then
      crc_var := crc_reg_8b;
      crc_err_8b <= '0';
      if TYPE_FRAME_DWI /= C_DATA_FRM then
        if end_CRC_8B_DWI = '1' then
          end_CRC_8B_DWI <= '0';
          if crc_reg_8b /= CRC_8B_DWI then
            crc_err_8b <= '1';
          end if;
          crc_reg_8b    <= (others => '0'); 

        elsif crc_to_inv_8b = '1' then
          crc_to_inv_8b <= '0';
          end_CRC_8B_DWI    <= '1'; 
          for i in 0 to 7 loop
            crc_var(i) := crc_reg_8b(7 - i); -- Bit-by-bit inversion
          end loop;
          crc_reg_8b <= crc_var; 

        elsif END_FRAME_DWI = '1'and NEW_WORD_DWI = '1'then
          crc_to_inv_8b <= '1';
          for i in indices_tier'range loop -- calculates the crc 8 byte by byte
              crc_var := calculate_crc_8(DATA_DWI(7+ indices_tier(i) downto 0 + indices_tier(i)), crc_var);
          end loop;
          crc_reg_8b <= crc_var; 

        elsif NEW_WORD_DWI = '1' then
          for i in indices'range loop -- calculates the crc 8 byte by byte
              crc_var := calculate_crc_8(DATA_DWI(7+ indices(i) downto 0 + indices(i)), crc_var);
          end loop;
          crc_reg_8b <= crc_var; 
        end if;
      end if;
    end if;
end process p_CRC_8B_DWI;

---------------------------------------------------------
-- Process: p_trans_ctrl_sig
-- Description: SEQ_NUM transmission
---------------------------------------------------------
p_trans_ctrl_sig: process(CLK, RST_N)
  variable crc_var : std_logic_vector(7 downto 0);
begin
  if RST_N = '0' then
    SEQ_NUM_DCCHECK    <= (others => '0'); 
    NEW_WORD_DCCHECK   <= '0'; 
    DATA_DCCHECK       <= (others => '0'); 
    TYPE_FRAME_DCCHECK <= (others => '0'); 
    CRC_ERR            <= '0';
    END_FRAME_DCCHECK  <= '0';
  elsif rising_edge(CLK) then
    SEQ_NUM_DCCHECK    <= SEQ_NUM_DWI;
    NEW_WORD_DCCHECK   <= NEW_WORD_DWI;
    END_FRAME_DCCHECK  <= END_FRAME_DWI;
    DATA_DCCHECK       <= DATA_DWI;
    TYPE_FRAME_DCCHECK <= TYPE_FRAME_DWI;
    if TYPE_FRAME_DWI = C_DATA_FRM then 
      CRC_ERR <= crc_err_16b;
    else
      CRC_ERR <= crc_err_8b;
    end if;
  end if;
end process p_trans_ctrl_sig;

end architecture rtl;