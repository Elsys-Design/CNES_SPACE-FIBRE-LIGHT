----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module describe the Data_word_id_fsm function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_word_id_fsm is
  port (
    RST_N                   : in  std_logic;                                    --! global reset
    CLK                     : in  std_logic;                                    --! Clock generated by GTY IP
    LINK_RESET              : in  std_logic;                                    --! Link Reset command 
    -- PHY PLUS LANE layer interface
    FIFO_RX_DATA_VALID_PPL  : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    FIFO_RX_RD_EN_PPL       : out  std_logic;                                   --! Flag to read data in FIFO RX  
    DATA_RX_PPL             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    VALID_K_CHARAC_PPL      : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);               --! K charachter valid in the 32-bit DATA_RX_PPL vector
    -- DCCHECK layer interface
    TYPE_FRAME_DWI          : out  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    NEW_WORD_DWI            : out  std_logic;   
    END_FRAME_DWI           : out  std_logic;
    DATA_DWI                : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    SEQ_NUM_DWI             : out  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX 
    CRC_16B_DWI             : out  std_logic_vector(15 downto 0);                --! Flag EMPTY of the FIFO RX
    CRC_8B_DWI              : out  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
    -- OTHER
    CRC_ERR                 : in   std_logic;   
    SEQ_ERR                 : in   std_logic;   
    FRAME_ERR               : out   std_logic;
		DETECTED_RXERR          : out std_logic  
  );
end data_word_id_fsm;

architecture rtl of data_word_id_fsm is

----------------------------- Declaration signals -----------------------------

-- Lane Initialisation FSM transition conditions process
   -- Type
type data_word_id_fsm_type is (
   RX_NOTHING_ST,                                                                --! Reset state
   RX_BROADCAST_FRAME_ST,                                                        --! Disabled TX and RX State
   RX_IDLE_FRAME_ST,                                                             --! Waiting State
   RX_DATA_FRAME_ST,                                                             --! Configuration INIT1 State
   RX_BROADCAST_AND_DATA_FRAME_ST
   );
   -- Signals
signal current_state                : data_word_id_fsm_type;                        --! Current state of the Dat Word Identification FSM
signal current_state_r              : data_word_id_fsm_type;                        --! Current state registered

signal receiving_frame    : std_logic;
signal type_incom_frame   : std_logic_vector(1 downto 0); 
signal data_word_cnt      : unsigned(7 downto 0); 
signal bc_word_cnt        : unsigned(1 downto 0);


signal detected_sdf     : std_logic ;
signal detected_edf     : std_logic ;
signal detected_sbf     : std_logic ;
signal detected_ebf     : std_logic ;
signal detected_sif     : std_logic ;
signal detected_fct     : std_logic ;
signal detected_ack     : std_logic ;
signal detected_nack    : std_logic ;
signal detected_full    : std_logic ;
signal detected_retry   : std_logic ;
signal detected_rxerr_i : std_logic ;

begin

	DETECTED_RXERR <= detected_rxerr_i;
-------------------------------------------------------------------------------------------
-- Data Word Identification FSM transition conditions process
p_fsm_data_word_id_transition : process(CLK,RST_N)
begin
   if RST_N = '0' then
      current_state     <= RX_NOTHING_ST;
      current_state_r   <= RX_NOTHING_ST;
      FRAME_ERR         <= '0';
   elsif rising_edge(CLK) then
      current_state_r   <= current_state;
      case current_state is
         when RX_NOTHING_ST                  => if LINK_RESET = '1' then
                                                   current_state  <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                   current_state  <= RX_BROADCAST_FRAME_ST;
                                                elsif detected_sdf ='1' then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_sif ='1' then
                                                   current_state  <= RX_IDLE_FRAME_ST;
                                                end if;
         when RX_DATA_FRAME_ST               => if LINK_RESET = '1' or detected_edf = '1' or detected_retry = '1' or detected_retry = '1' or CRC_ERR = '1' or SEQ_ERR = '1' then
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif detected_sdf = '1' or detected_sif = '1' or detected_ebf = '1' or data_word_cnt > C_MAX_DATA_FRAME then
                                                  FRAME_ERR      <= '1';
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                  current_state  <= RX_BROADCAST_AND_DATA_FRAME_ST;
                                                end if;
         when RX_BROADCAST_FRAME_ST          => if LINK_RESET = '1' or (detected_ebf = '1' and bc_word_cnt = C_WORD_BC_FRAME) or detected_retry = '1' or detected_retry = '1' or CRC_ERR = '1' or SEQ_ERR = '1' then
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif detected_sdf = '1' or detected_sbf = '1' or detected_sif = '1' or detected_edf = '1' or (detected_ebf = '1' and bc_word_cnt /= C_WORD_BC_FRAME) or bc_word_cnt > C_WORD_BC_FRAME then
                                                   FRAME_ERR      <= '1';
                                                   current_state  <= RX_NOTHING_ST;
                                                end if;
      
         when RX_BROADCAST_AND_DATA_FRAME_ST => if LINK_RESET = '1' or detected_retry = '1' or detected_retry = '1' or CRC_ERR = '1' or SEQ_ERR = '1' then
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif (detected_ebf = '1' and bc_word_cnt = C_WORD_BC_FRAME) then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_sdf = '1' or detected_sbf = '1' or detected_sif = '1' or detected_edf = '1' or (detected_ebf = '1' and bc_word_cnt /= C_WORD_BC_FRAME) or bc_word_cnt > C_WORD_BC_FRAME then
                                                   FRAME_ERR      <= '1';
                                                   current_state  <= RX_NOTHING_ST;
                                                end if;
      
         when RX_IDLE_FRAME_ST               => if LINK_RESET = '1' or detected_retry = '1' or detected_retry = '1' or CRC_ERR = '1' or SEQ_ERR = '1' then
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                   current_state  <= RX_BROADCAST_FRAME_ST;
                                                elsif detected_sdf ='1' then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_edf = '1' or detected_ebf = '1' or data_word_cnt > C_MAX_IDLE_FRAME then
                                                   FRAME_ERR      <= '1';
                                                   current_state  <= RX_NOTHING_ST;
                                                end if;
         when others                          => current_state  <= RX_NOTHING_ST;
      end case;
   end if;
end process p_fsm_data_word_id_transition;

-- Data Word Identification FSM action on state process
p_comb_state : process(CLK,RST_N)
begin
	if RST_N = '0' then
	   receiving_frame         <= '0';
	   type_incom_frame        <= (others =>'0');
	   data_word_cnt           <= (others =>'0');
	   bc_word_cnt             <= (others =>'0');
	elsif rising_edge(CLK) then
		if current_state = RX_NOTHING_ST then
		  receiving_frame      <= '0';
		  data_word_cnt        <= (others =>'0');
		  bc_word_cnt          <= (others =>'0');
		elsif current_state = RX_DATA_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "01";               -- receiving data frame
		  if (current_state_r = RX_IDLE_FRAME_ST) then
		    data_word_cnt      <= to_unsigned(1,data_word_cnt'length);
		  else
		    data_word_cnt      <= data_word_cnt + 1;
		  end if; 
		elsif current_state = RX_BROADCAST_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "10";               -- receiving broadcast frame
		  bc_word_cnt          <= bc_word_cnt + 1;
		  data_word_cnt        <= (others =>'0');
		elsif current_state = RX_BROADCAST_AND_DATA_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "10";               -- receiving broadcast frame
		  bc_word_cnt          <= bc_word_cnt + 1;
		elsif current_state = RX_IDLE_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "11";               -- receiving idle frame
		  data_word_cnt        <= data_word_cnt + 1;
		end if;
	end if;
end process p_comb_state;

-- Data Word Identification FSM action on state process
p_data_word_detection : process(CLK,RST_N)
begin
	if RST_N = '0' then
		detected_sdf     <= '0';
		NEW_WORD_DWI     <= '0';
		detected_edf     <= '0';
		detected_sbf     <= '0';
		detected_ebf     <= '0';
		detected_sif     <= '0';
		detected_fct     <= '0';
		detected_ack     <= '0';
		detected_nack    <= '0';
		detected_full    <= '0';
		detected_retry   <= '0';
		detected_rxerr_i   <= '0';
    SEQ_NUM_DWI      <= (others=> '0');
    CRC_16B_DWI      <= (others=> '0');
    CRC_8B_DWI       <= (others=> '0');
		TYPE_FRAME_DWI   <= (others=> '0');
		DATA_DWI         <= (others=> '0');
    END_FRAME_DWI    <= '0';
	elsif rising_edge(CLK) then
		-- Reset of signals
		detected_sdf     <= '0';
		detected_edf     <= '0';
		detected_sbf     <= '0';
		detected_ebf     <= '0';
		detected_sif     <= '0';
		detected_fct     <= '0';
		detected_ack     <= '0';
		detected_nack    <= '0';
		detected_full    <= '0';
		detected_retry   <= '0';
		detected_rxerr_i   <= '0';
    END_FRAME_DWI    <= '0';
		-- Frame treatment
	  if (FIFO_RX_DATA_VALID_PPL ='1') then 
			if current_state = RX_IDLE_FRAME_ST then
				DATA_DWI       <= DATA_RX_PPL;
        NEW_WORD_DWI   <= '0';
	  	elsif DATA_RX_PPL(15 downto 0) = C_SDF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SDF control word detected
	  		detected_sdf   <= '1';                                                -- Set SDF flag detected to '1'
	  		TYPE_FRAME_DWI <= C_DATA_FRM;
	  		NEW_WORD_DWI   <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_0_SYMB and VALID_K_CHARAC_PPL = "0001" then -- EDF control word detected
	  		detected_edf   <= '1'; 
	  		TYPE_FRAME_DWI <= C_DATA_FRM;                                                   -- Set EDF flag detected to '1'
	  		NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    <= DATA_RX_PPL(15 downto 8);
	  		CRC_16B_DWI    <= DATA_RX_PPL(31 downto 16); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_SBF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SBF control word detected
	  		detected_sbf   <= '1'; 
	  		TYPE_FRAME_DWI <= C_BC_FRM;                                                  -- Set SBF flag detected to '1'
	  		NEW_WORD_DWI   <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_2_SYMB and VALID_K_CHARAC_PPL = "0001" then -- EBF control word detected
	  		detected_ebf   <= '1';                                                    -- Set EBF flag detected to '1'
	  		TYPE_FRAME_DWI <= C_BC_FRM;   
	  		NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16); 
	  		CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_SIF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SIF control word detected
	  		detected_sif   <= '1';                                                   -- Set SIF flag detected to '1'
	  		TYPE_FRAME_DWI <= C_IDLE_FRM;   
	  		NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16); 
	  		CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_3_SYMB and VALID_K_CHARAC_PPL = "0001" then -- FCT control word detected
	  		detected_fct   <= '1';                                                    -- Set FCT flag detected to '1'
	  		TYPE_FRAME_DWI <= C_FCT_FRM; 
	  		NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16);
	  		CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_ACK_WORD and VALID_K_CHARAC_PPL = "0001" then -- ACK control word detected
	  	  detected_ack   <= '1';                                                   -- Set ACK flag detected to '1'
	  	  TYPE_FRAME_DWI <= C_ACK_FRM;
	  	  NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_NACK_WORD and VALID_K_CHARAC_PPL = "0001" then -- NACK control word detected
	  	  detected_nack  <= '1';                                                    -- Set NACK flag detected to '1'
	  	  TYPE_FRAME_DWI <= C_NACK_FRM;
	  	  NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_FULL_WORD and VALID_K_CHARAC_PPL = "0001" then -- FULL control word detected
	  	  detected_full  <= '1';                                                    -- Set FULL flag detected to '1'
	  	  TYPE_FRAME_DWI <= C_FULL_FRM;
	  	  NEW_WORD_DWI   <= '1';
        END_FRAME_DWI  <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL(15 downto 0) = C_RETRY_WORD and VALID_K_CHARAC_PPL = "0001" then -- RETRY control word detected
	  	  detected_retry <= '1';                                                     -- Set RETRY flag detected to '1'
	  	  TYPE_FRAME_DWI <= C_RETRY_FRM;
	  	  NEW_WORD_DWI   <= '1';
				DATA_DWI       <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     <= DATA_RX_PPL(31 downto 24); 
	  	elsif DATA_RX_PPL = C_RXERR_WORD and VALID_K_CHARAC_PPL = "0001" then -- RXERR control word detected
	  	  detected_rxerr_i <= '1';                                         -- Set RXERR flag detected to '1'
        NEW_WORD_DWI   <= '0';
      else
        DATA_DWI       <= DATA_RX_PPL;
        NEW_WORD_DWI   <= '1';
	  	end if;
    else
      NEW_WORD_DWI     <= '0';
	  end if;
	end if;
end process p_data_word_detection;

---------------------------------------------------------
-- Process: p_fifo_rd_ppl
-- Description: Write frames into the fifo
---------------------------------------------------------
p_fifo_rd_ppl: process(CLK, RST_N)
begin
	if RST_N = '0' then
		FIFO_RX_RD_EN_PPL <= '0';
	elsif rising_edge(CLK) then
		FIFO_RX_RD_EN_PPL <= '1';
	end if;
end process p_fifo_rd_ppl;  

end architecture rtl;