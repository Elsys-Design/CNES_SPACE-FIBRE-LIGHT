-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 23/07/2025
--
-- Description : This is the testbench of the ppl_64_lane_ctrl_word_detect module
----------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library work;
   use work.pkg_simu.all;

entity tb_ppl_64_lane_ctrl_word_detect is
end entity;

architecture tb of tb_ppl_64_lane_ctrl_word_detect is

component ppl_64_lane_ctrl_word_detect is
  port (
    RST_N                            : in  std_logic;                                    --! Global reset. Active Low
    CLK                              : in  std_logic;                                    --! Clock generated by HSSL IP
    -- ppl_64_lane_init_fsm (PLIF) interface
    NO_SIGNAL_PLCWD                  : out std_logic;                                    --! Flag indicating that no signal is received
    RX_NEW_WORD_PLCWD                : out std_logic_vector(1 downto 0);                 --! Flag indicating that a new word has been received
    DETECTED_INIT1_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT1 control word received
    DETECTED_INIT2_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT2 control word received
    DETECTED_INIT3_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT3 control word received
    DETECTED_INV_INIT1_PLCWD         : out std_logic_vector(1 downto 0);                 --! Flag indicating INV_INIT1 control word received
    DETECTED_INV_INIT2_PLCWD         : out std_logic_vector(1 downto 0);                 --! Flag indicating INV_INIT2 control word received
    DETECTED_RXERR_WORD_PLCWD        : out std_logic_vector(1 downto 0);                 --! Flag indicating RXERR control word detected
    DETECTED_LOSS_SIGNAL_PLCWD       : out std_logic_vector(1 downto 0);                 --! Flag indicating LOSS_SIGNAL control word detected
    DETECTED_STANDBY_PLCWD           : out std_logic_vector(1 downto 0);                 --! Flag indicating STANDBY control word detected
    COMMA_K287_RXED_PLCWD            : out std_logic_vector(1 downto 0);                 --! Comma K28.7 character received flag
    CAPABILITY_PLCWD                 : out std_logic_vector(15 downto 0);                --! Capability extracted from INIT3 control word: bits [31:24] and [63:56]
    SEND_RXERR_PLIF                  : in  std_logic_vector(1 downto 0);                 --! Flag to send RXERR control word to Data-Link layer when FSM exits ACTIVE_ST
    NO_SIGNAL_DETECTION_ENABLED_PLIF : in  std_logic;                                    --! Flag to enable the no-signal detection function
    ENABLE_TRANSM_DATA_PLIF          : in  std_logic;                                    --! Flag to enable the transmission of data
    -- ppl_64_parallel_loopback (PLPL) interface
    DATA_RX_PLPL                     : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data from ppl_64_parallel_loopback
    VALID_K_CHARAC_PLPL              : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags from ppl_64_parallel_loopback
    DATA_RDY_PLPL                    : in  std_logic;                                    --! Data valid flag from ppl_64_parallel_loopback
    LOSS_OF_SIGNAL_PLPL              : in  std_logic;                                    --! Loss of signal flag from ppl_64_parallel_loopback
    -- ppl_64_rx_wr_en_fifo (PLRWEF) interface
    DATA_RX_PLCWD                    : out std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data sent to Data-Link layer
    VALID_K_CHARAC_PLCWD             : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags sent to Data-Link layer
    DATA_RDY_PLCWD                   : out std_logic_vector(1 downto 0)                  --! Data valid flag sent to Data-Link layer
  );
end component;


---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
constant periode                        : time := 13.334 ns;

signal RST_N                            : std_logic := '0';
signal CLK                              : std_logic := '0';

signal NO_SIGNAL_PLCWD                  : std_logic;
signal RX_NEW_WORD_PLCWD                : std_logic_vector(1 downto 0);
signal DETECTED_INIT1_PLCWD             : std_logic_vector(1 downto 0);
signal DETECTED_INIT2_PLCWD             : std_logic_vector(1 downto 0);
signal DETECTED_INIT3_PLCWD             : std_logic_vector(1 downto 0);
signal DETECTED_INV_INIT1_PLCWD         : std_logic_vector(1 downto 0);
signal DETECTED_INV_INIT2_PLCWD         : std_logic_vector(1 downto 0);
signal DETECTED_RXERR_WORD_PLCWD        : std_logic_vector(1 downto 0);
signal DETECTED_LOSS_SIGNAL_PLCWD       : std_logic_vector(1 downto 0);
signal DETECTED_STANDBY_PLCWD           : std_logic_vector(1 downto 0);
signal COMMA_K287_RXED_PLCWD            : std_logic_vector(1 downto 0);
signal CAPABILITY_PLCWD                 : std_logic_vector(15 downto 0);
signal SEND_RXERR_PLIF                  : std_logic_vector(1 downto 0) := "00";
signal NO_SIGNAL_DETECTION_ENABLED_PLIF : std_logic := '0';
signal ENABLE_TRANSM_DATA_PLIF          : std_logic := '0';
signal DATA_RX_PLPL                     : std_logic_vector(C_DATA_WIDTH-1 downto 0)  := (others =>'0');
signal VALID_K_CHARAC_PLPL              : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0):= (others =>'0');
signal DATA_RDY_PLPL                    : std_logic := '0';
signal LOSS_OF_SIGNAL_PLPL              : std_logic := '1';
signal DATA_RX_PLCWD                    : std_logic_vector(C_DATA_WIDTH-1 downto 0);
signal VALID_K_CHARAC_PLCWD             : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
signal DATA_RDY_PLCWD                   : std_logic_vector(1 downto 0);

signal capability_in                    : std_logic_vector(7 downto 0):= (others => '0');
signal lost_cause                       : std_logic_vector(1 downto 0):= (others => '0');
signal standby_reason                   : std_logic_vector(7 downto 0):= (others => '0');
begin

---------------------------------------------------------
-----                  Instantiation                -----
---------------------------------------------------------
DUT : ppl_64_lane_ctrl_word_detect
port map(
  RST_N                            => RST_N,
  CLK                              => CLK,
  NO_SIGNAL_PLCWD                  => NO_SIGNAL_PLCWD,
  RX_NEW_WORD_PLCWD                => RX_NEW_WORD_PLCWD,
  DETECTED_INIT1_PLCWD             => DETECTED_INIT1_PLCWD,
  DETECTED_INIT2_PLCWD             => DETECTED_INIT2_PLCWD,
  DETECTED_INIT3_PLCWD             => DETECTED_INIT3_PLCWD,
  DETECTED_INV_INIT1_PLCWD         => DETECTED_INV_INIT1_PLCWD,
  DETECTED_INV_INIT2_PLCWD         => DETECTED_INV_INIT2_PLCWD,
  DETECTED_RXERR_WORD_PLCWD        => DETECTED_RXERR_WORD_PLCWD,
  DETECTED_LOSS_SIGNAL_PLCWD       => DETECTED_LOSS_SIGNAL_PLCWD,
  DETECTED_STANDBY_PLCWD           => DETECTED_STANDBY_PLCWD,
  COMMA_K287_RXED_PLCWD            => COMMA_K287_RXED_PLCWD,
  CAPABILITY_PLCWD                 => CAPABILITY_PLCWD,
  SEND_RXERR_PLIF                  => SEND_RXERR_PLIF,
  NO_SIGNAL_DETECTION_ENABLED_PLIF => NO_SIGNAL_DETECTION_ENABLED_PLIF,
  ENABLE_TRANSM_DATA_PLIF          => ENABLE_TRANSM_DATA_PLIF,
  DATA_RX_PLPL                     => DATA_RX_PLPL,
  VALID_K_CHARAC_PLPL              => VALID_K_CHARAC_PLPL,
  DATA_RDY_PLPL                    => DATA_RDY_PLPL,
  LOSS_OF_SIGNAL_PLPL              => LOSS_OF_SIGNAL_PLPL,
  DATA_RX_PLCWD                    => DATA_RX_PLCWD,
  VALID_K_CHARAC_PLCWD             => VALID_K_CHARAC_PLCWD,
  DATA_RDY_PLCWD                   => DATA_RDY_PLCWD
);

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
-- generate clock 150 MHz
horloge : process
begin
   CLK   <= not CLK;
   wait for periode/2;
end process;

scenario : process
  variable test_failed : boolean := false;
begin
  RST_N <= '0';
  wait for 10 us;
  wait until rising_edge(CLK);
  RST_N <= '1';
  wait for 20 us;
  DATA_RDY_PLPL           <= '1';
  ENABLE_TRANSM_DATA_PLIF <= '1';
  wait for 1 us;
  capability_in      <= x"FF";
  lost_cause         <= "11";
  standby_reason     <= x"DD";
  wait until rising_edge(CLK);
  wait until falling_edge(CLK);
  --------------------------------------
  -- TEST 0: INIT1 detect             --
  --------------------------------------
  -- Test 0.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_INIT1_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 0.1: INIT 1: DATA_RX_PLCWD",        x"12345678"& x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 0.1: INIT 1: VALID_K_CHARAC_PLCWD", x"00",                    VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 0.1: INIT 1: DATA_RDY_PLCWD",       "10",                     DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 0.1: INIT 1: RX_NEW_WORD_PLCWD",    "11",                     RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 0.1: INIT 1: DETECTED_INIT1_PLCWD", "01",                     DETECTED_INIT1_PLCWD, test_failed);

  -- Test 0.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_INIT1_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 0.2: INIT 1: DATA_RX_PLCWD",        x"00000000" & x"12345678", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 0.2: INIT 1: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 0.2: INIT 1: DATA_RDY_PLCWD",       "01",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 0.2: INIT 1: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 0.2: INIT 1: DETECTED_INIT1_PLCWD", "10",                      DETECTED_INIT1_PLCWD, test_failed);

  -- Test 0.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_INIT1_WORD & C_INIT1_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 0.3: INIT 1: DATA_RX_PLCWD",        x"00000000" & x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 0.3: INIT 1: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 0.3: INIT 1: DATA_RDY_PLCWD",       "00",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 0.3: INIT 1: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 0.3: INIT 1: DETECTED_INIT1_PLCWD", "11",                      DETECTED_INIT1_PLCWD, test_failed);

  --------------------------------------
  -- TEST 1: INIT2 detect             --
  --------------------------------------
  -- Test 1.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_INIT2_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 1.1: INIT 2: DATA_RX_PLCWD",        x"12345678"& x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 1.1: INIT 2: VALID_K_CHARAC_PLCWD", x"00",                    VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 1.1: INIT 2: DATA_RDY_PLCWD",       "10",                     DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 1.1: INIT 2: RX_NEW_WORD_PLCWD",    "11",                     RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 1.1: INIT 2: DETECTED_INIT2_PLCWD", "01",                     DETECTED_INIT2_PLCWD, test_failed);

  -- Test 1.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_INIT2_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 1.2: INIT 2: DATA_RX_PLCWD",        x"00000000" & x"12345678", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 1.2: INIT 2: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 1.2: INIT 2: DATA_RDY_PLCWD",       "01",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 1.2: INIT 2: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 1.2: INIT 2: DETECTED_INIT2_PLCWD", "10",                      DETECTED_INIT2_PLCWD, test_failed);

  -- Test 1.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_INIT2_WORD & C_INIT2_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 1.3: INIT 2: DATA_RX_PLCWD",        x"00000000" & x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 1.3: INIT 2: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 1.3: INIT 2: DATA_RDY_PLCWD",       "00",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 1.3: INIT 2: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 1.3: INIT 2: DETECTED_INIT2_PLCWD", "11",                      DETECTED_INIT2_PLCWD, test_failed);

  --------------------------------------
  -- TEST 2: INIT3 detect             --
  --------------------------------------
  -- Test 2.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& capability_in & C_INIT3_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 2.1: INIT 3: DATA_RX_PLCWD",        x"12345678"& x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 2.1: INIT 3: CAPABILITY_PLCWD",     x"00" & x"FF",            CAPABILITY_PLCWD,     test_failed);
  check_equal("Test 2.1: INIT 3: VALID_K_CHARAC_PLCWD", x"00",                    VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 2.1: INIT 3: DATA_RDY_PLCWD",       "10",                     DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 2.1: INIT 3: RX_NEW_WORD_PLCWD",    "11",                     RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 2.1: INIT 3: DETECTED_INIT3_PLCWD", "01",                     DETECTED_INIT3_PLCWD, test_failed);

  -- Test 2.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= capability_in & C_INIT3_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 2.2: INIT 3: DATA_RX_PLCWD",        x"00000000" & x"12345678", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 2.2: INIT 3: CAPABILITY_PLCWD",     x"FF" & x"00",             CAPABILITY_PLCWD,     test_failed);
  check_equal("Test 2.2: INIT 3: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 2.2: INIT 3: DATA_RDY_PLCWD",       "01",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 2.2: INIT 3: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 2.2: INIT 3: DETECTED_INIT3_PLCWD", "10",                      DETECTED_INIT3_PLCWD, test_failed);

  -- Test 2.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= capability_in & C_INIT3_WORD & capability_in & C_INIT3_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 2.3: INIT 3: DATA_RX_PLCWD",        x"00000000" & x"00000000", DATA_RX_PLCWD,        test_failed);
  check_equal("Test 2.3: INIT 3: CAPABILITY_PLCWD",     x"FF" & x"FF",             CAPABILITY_PLCWD,     test_failed);
  check_equal("Test 2.3: INIT 3: VALID_K_CHARAC_PLCWD", x"00",                     VALID_K_CHARAC_PLCWD, test_failed);
  check_equal("Test 2.3: INIT 3: DATA_RDY_PLCWD",       "00",                      DATA_RDY_PLCWD,       test_failed);
  check_equal("Test 2.3: INIT 3: RX_NEW_WORD_PLCWD",    "11",                      RX_NEW_WORD_PLCWD,    test_failed);
  check_equal("Test 2.3: INIT 3: DETECTED_INIT3_PLCWD", "11",                      DETECTED_INIT3_PLCWD, test_failed);

  --------------------------------------
  -- TEST 3: iINIT1 detect             --
  --------------------------------------
  -- Test 3.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_I_INIT1_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 3.1: iINIT 1: DATA_RX_PLCWD",            x"12345678"& x"00000000", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 3.1: iINIT 1: VALID_K_CHARAC_PLCWD",     x"00",                    VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 3.1: iINIT 1: DATA_RDY_PLCWD",           "10",                     DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 3.1: iINIT 1: RX_NEW_WORD_PLCWD",        "11",                     RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 3.1: iINIT 1: DETECTED_INV_INIT1_PLCWD", "01",                     DETECTED_INV_INIT1_PLCWD, test_failed);

  -- Test 3.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_I_INIT1_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 3.2: iINIT 1: DATA_RX_PLCWD",            x"00000000" & x"12345678", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 3.2: iINIT 1: VALID_K_CHARAC_PLCWD",     x"00",                     VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 3.2: iINIT 1: DATA_RDY_PLCWD",           "01",                      DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 3.2: iINIT 1: RX_NEW_WORD_PLCWD",        "11",                      RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 3.2: iINIT 1: DETECTED_INV_INIT1_PLCWD", "10",                      DETECTED_INV_INIT1_PLCWD, test_failed);

  -- Test 3.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_I_INIT1_WORD & C_I_INIT1_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 3.3: iINIT 1: DATA_RX_PLCWD",            x"00000000" & x"00000000", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 3.3: iINIT 1: VALID_K_CHARAC_PLCWD",     x"00",                     VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 3.3: iINIT 1: DATA_RDY_PLCWD",           "00",                      DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 3.3: iINIT 1: RX_NEW_WORD_PLCWD",        "11",                      RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 3.3: iINIT 1: DETECTED_INV_INIT1_PLCWD", "11",                      DETECTED_INV_INIT1_PLCWD, test_failed);

  --------------------------------------
  -- TEST 4: iINIT2 detect             --
  --------------------------------------
  -- Test 4.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_I_INIT2_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 4.1: iINIT 2: DATA_RX_PLCWD",            x"12345678"& x"00000000", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 4.1: iINIT 2: VALID_K_CHARAC_PLCWD",     x"00",                    VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 4.1: iINIT 2: DATA_RDY_PLCWD",           "10",                     DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 4.1: iINIT 2: RX_NEW_WORD_PLCWD",        "11",                     RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 4.1: iINIT 2: DETECTED_INV_INIT2_PLCWD", "01",                     DETECTED_INV_INIT2_PLCWD, test_failed);

  -- Test 4.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_I_INIT2_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 4.2: iINIT 2: DATA_RX_PLCWD",            x"00000000" & x"12345678", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 4.2: iINIT 2: VALID_K_CHARAC_PLCWD",     x"00",                     VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 4.2: iINIT 2: DATA_RDY_PLCWD",           "01",                      DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 4.2: iINIT 2: RX_NEW_WORD_PLCWD",        "11",                      RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 4.2: iINIT 2: DETECTED_INV_INIT2_PLCWD", "10",                      DETECTED_INV_INIT2_PLCWD, test_failed);

  -- Test 4.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_I_INIT2_WORD & C_I_INIT2_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 4.3: iINIT 2: DATA_RX_PLCWD",            x"00000000" & x"00000000", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 4.3: iINIT 2: VALID_K_CHARAC_PLCWD",     x"00",                     VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 4.3: iINIT 2: DATA_RDY_PLCWD",           "00",                      DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 4.3: iINIT 2: RX_NEW_WORD_PLCWD",        "11",                      RX_NEW_WORD_PLCWD,        test_failed);
  check_equal("Test 4.3: iINIT 2: DETECTED_INV_INIT2_PLCWD", "11",                      DETECTED_INV_INIT2_PLCWD, test_failed);

  --------------------------------------
  -- TEST 5: LOST SIGNAL detect       --
  --------------------------------------
  -- Test 5.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& "000000" & lost_cause & C_LOST_SIG_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 5.1: LOST SIGNAL: DATA_RX_PLCWD",              x"12345678"& x"00000000", DATA_RX_PLCWD,              test_failed);
  check_equal("Test 5.1: LOST SIGNAL: COMMA_K287_RXED_PLCWD",      "01",                     COMMA_K287_RXED_PLCWD,      test_failed);
  check_equal("Test 5.1: LOST SIGNAL: VALID_K_CHARAC_PLCWD",       x"00",                    VALID_K_CHARAC_PLCWD,       test_failed);
  check_equal("Test 5.1: LOST SIGNAL: DATA_RDY_PLCWD",             "10",                     DATA_RDY_PLCWD,             test_failed);
  check_equal("Test 5.1: LOST SIGNAL: RX_NEW_WORD_PLCWD",          "11",                     RX_NEW_WORD_PLCWD,          test_failed);
  check_equal("Test 5.1: LOST SIGNAL: DETECTED_LOSS_SIGNAL_PLCWD", "01",                     DETECTED_LOSS_SIGNAL_PLCWD, test_failed);

  -- Test 5.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= "000000" & lost_cause & C_LOST_SIG_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 5.2: LOST SIGNAL: DATA_RX_PLCWD",              x"00000000" & x"12345678", DATA_RX_PLCWD,              test_failed);
  check_equal("Test 5.2: LOST SIGNAL: COMMA_K287_RXED_PLCWD",      "10",                      COMMA_K287_RXED_PLCWD,      test_failed);
  check_equal("Test 5.2: LOST SIGNAL: VALID_K_CHARAC_PLCWD",       x"00",                     VALID_K_CHARAC_PLCWD,       test_failed);
  check_equal("Test 5.2: LOST SIGNAL: DATA_RDY_PLCWD",             "01",                      DATA_RDY_PLCWD,             test_failed);
  check_equal("Test 5.2: LOST SIGNAL: RX_NEW_WORD_PLCWD",          "11",                      RX_NEW_WORD_PLCWD,          test_failed);
  check_equal("Test 5.2: LOST SIGNAL: DETECTED_LOSS_SIGNAL_PLCWD", "10",                      DETECTED_LOSS_SIGNAL_PLCWD, test_failed);

  -- Test 5.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= "000000" & lost_cause & C_LOST_SIG_WORD & "000000" & lost_cause & C_LOST_SIG_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 5.3: LOST SIGNAL: DATA_RX_PLCWD",              x"00000000" & x"00000000", DATA_RX_PLCWD,              test_failed);
  check_equal("Test 5.3: LOST SIGNAL: COMMA_K287_RXED_PLCWD",      "11" ,                     COMMA_K287_RXED_PLCWD,      test_failed);
  check_equal("Test 5.3: LOST SIGNAL: VALID_K_CHARAC_PLCWD",       x"00",                     VALID_K_CHARAC_PLCWD,       test_failed);
  check_equal("Test 5.3: LOST SIGNAL: DATA_RDY_PLCWD",             "00",                      DATA_RDY_PLCWD,             test_failed);
  check_equal("Test 5.3: LOST SIGNAL: RX_NEW_WORD_PLCWD",          "11",                      RX_NEW_WORD_PLCWD,          test_failed);
  check_equal("Test 5.3: LOST SIGNAL: DETECTED_LOSS_SIGNAL_PLCWD", "11",                      DETECTED_LOSS_SIGNAL_PLCWD, test_failed);

  --------------------------------------
  -- TEST 6: STANDBY detect       --
  --------------------------------------
  -- Test 6.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& standby_reason & C_STANDBY_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 6.1: STANDBY: DATA_RX_PLCWD",          x"12345678"& x"00000000", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 6.1: STANDBY: COMMA_K287_RXED_PLCWD",  "01",                     COMMA_K287_RXED_PLCWD,  test_failed);
  check_equal("Test 6.1: STANDBY: VALID_K_CHARAC_PLCWD",   x"00",                    VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 6.1: STANDBY: DATA_RDY_PLCWD",         "10",                     DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 6.1: STANDBY: RX_NEW_WORD_PLCWD",      "11",                     RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 6.1: STANDBY: DETECTED_STANDBY_PLCWD", "01",                     DETECTED_STANDBY_PLCWD, test_failed);

  -- Test 6.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= standby_reason & C_STANDBY_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 6.2: STANDBY: DATA_RX_PLCWD",          x"00000000" & x"12345678", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 6.2: STANDBY: COMMA_K287_RXED_PLCWD",  "10",                      COMMA_K287_RXED_PLCWD,  test_failed);
  check_equal("Test 6.2: STANDBY: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 6.2: STANDBY: DATA_RDY_PLCWD",         "01",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 6.2: STANDBY: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 6.2: STANDBY: DETECTED_STANDBY_PLCWD", "10",                      DETECTED_STANDBY_PLCWD, test_failed);

  -- Test 6.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= standby_reason & C_STANDBY_WORD & standby_reason & C_STANDBY_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 6.3: STANDBY: DATA_RX_PLCWD",          x"00000000" & x"00000000", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 6.3: STANDBY: COMMA_K287_RXED_PLCWD",  "11",                      COMMA_K287_RXED_PLCWD,  test_failed);
  check_equal("Test 6.3: STANDBY: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 6.3: STANDBY: DATA_RDY_PLCWD",         "00",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 6.3: STANDBY: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 6.3: STANDBY: DETECTED_STANDBY_PLCWD", "11",                      DETECTED_STANDBY_PLCWD, test_failed);

  --------------------------------------
  -- TEST 7: Send RXERR detect        --
  --------------------------------------
  -- Test 7.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678" & x"12345678";
  VALID_K_CHARAC_PLPL <= x"0" & x"0";
  SEND_RXERR_PLIF    <= "01";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 7.1: RXERR: DATA_RX_PLCWD",            x"12345678" & C_RXERR_WORD, DATA_RX_PLCWD,            test_failed);
  check_equal("Test 7.1: RXERR: VALID_K_CHARAC_PLCWD",     x"01",                      VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 7.1: RXERR: DATA_RDY_PLCWD",           "11",                       DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 7.1: RXERR: RX_NEW_WORD_PLCWD",        "10",                       RX_NEW_WORD_PLCWD,        test_failed);

  -- Test 7.2: Second word only
  --------------------------------------
  SEND_RXERR_PLIF    <= "10";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 7.2: RXERR: DATA_RX_PLCWD",            C_RXERR_WORD & x"12345678", DATA_RX_PLCWD,            test_failed);
  check_equal("Test 7.2: RXERR: VALID_K_CHARAC_PLCWD",     x"10",                      VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 7.2: RXERR: DATA_RDY_PLCWD",           "11",                       DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 7.2: RXERR: RX_NEW_WORD_PLCWD",        "01",                       RX_NEW_WORD_PLCWD,        test_failed);

  -- Test 7.3: 2 words
  --------------------------------------
  SEND_RXERR_PLIF    <= "11";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 7.3: RXERR: DATA_RX_PLCWD",            C_RXERR_WORD & C_RXERR_WORD, DATA_RX_PLCWD,            test_failed);
  check_equal("Test 7.3: RXERR: VALID_K_CHARAC_PLCWD",     x"11",                       VALID_K_CHARAC_PLCWD,     test_failed);
  check_equal("Test 7.3: RXERR: DATA_RDY_PLCWD",           "11",                        DATA_RDY_PLCWD,           test_failed);
  check_equal("Test 7.3: RXERR: RX_NEW_WORD_PLCWD",        "00",                        RX_NEW_WORD_PLCWD,        test_failed);
  SEND_RXERR_PLIF    <= "00";
  --------------------------------------
  -- TEST 8: Transmit DATA            --
  --------------------------------------
  -- Test 8.1: 2 data words
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678" & x"9abcdef0";
  VALID_K_CHARAC_PLPL <= x"0" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 8.1: DATA: DATA_RX_PLCWD",             x"12345678" & x"9abcdef0", DATA_RX_PLCWD,             test_failed);
  check_equal("Test 8.1: DATA: VALID_K_CHARAC_PLCWD",      x"00",                     VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 8.1: DATA: DATA_RDY_PLCWD",            "11",                      DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 8.1: DATA: RX_NEW_WORD_PLCWD",         "11",                      RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 8.1: DATA: DETECTED_RXERR_WORD_PLCWD", "00",                      DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 8.2: First word only RXERR
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678" & C_RXERR_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 8.2: DATA: DATA_RX_PLCWD",             x"12345678" & C_RXERR_WORD, DATA_RX_PLCWD,             test_failed);
  check_equal("Test 8.2: DATA: VALID_K_CHARAC_PLCWD",      x"01",                      VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 8.2: DATA: DATA_RDY_PLCWD",            "11",                       DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 8.2: DATA: RX_NEW_WORD_PLCWD",         "11",                       RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 8.2: DATA: DETECTED_RXERR_WORD_PLCWD", "01",                       DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 8.3: Second word only RXERR
  --------------------------------------
  DATA_RX_PLPL       <= C_RXERR_WORD & x"9abcdef0";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 8.3: DATA: DATA_RX_PLCWD",             C_RXERR_WORD & x"9abcdef0", DATA_RX_PLCWD,             test_failed);
  check_equal("Test 8.3: DATA: VALID_K_CHARAC_PLCWD",      x"10",                      VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 8.3: DATA: DATA_RDY_PLCWD",            "11",                       DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 8.3: DATA: RX_NEW_WORD_PLCWD",         "11",                       RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 8.1: DATA: DETECTED_RXERR_WORD_PLCWD", "10",                       DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 8.4: 2 words RXERR
  --------------------------------------
  DATA_RX_PLPL       <= C_RXERR_WORD & C_RXERR_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 8.4: DATA: DATA_RX_PLCWD",             C_RXERR_WORD & C_RXERR_WORD, DATA_RX_PLCWD,             test_failed);
  check_equal("Test 8.4: DATA: VALID_K_CHARAC_PLCWD",      x"11",                       VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 8.4: DATA: DATA_RDY_PLCWD",            "11",                        DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 8.4: DATA: RX_NEW_WORD_PLCWD",         "11",                        RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 8.4: DATA: DETECTED_RXERR_WORD_PLCWD", "11",                        DETECTED_RXERR_WORD_PLCWD, test_failed);

  --------------------------------------
  -- TEST 9: SKIP detect             --
  --------------------------------------
  -- Test 9.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_SKIP_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 9.1: SKIP: DATA_RX_PLCWD",          x"12345678"& x"00000000", DATA_RX_PLCWD,           test_failed);
  check_equal("Test 9.1: SKIP: VALID_K_CHARAC_PLCWD",   x"00",                    VALID_K_CHARAC_PLCWD,    test_failed);
  check_equal("Test 9.1: SKIP: DATA_RDY_PLCWD",         "10",                     DATA_RDY_PLCWD,          test_failed);
  check_equal("Test 9.1: SKIP: RX_NEW_WORD_PLCWD",      "11",                     RX_NEW_WORD_PLCWD,       test_failed);
  check_equal("Test 9.1: SKIP: COMMA_K287_RXED_PLCWD",  "01",                     COMMA_K287_RXED_PLCWD,   test_failed);

  -- Test 9.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_SKIP_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 9.2: SKIP: DATA_RX_PLCWD",          x"00000000" & x"12345678", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 9.2: SKIP: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 9.2: SKIP: DATA_RDY_PLCWD",         "01",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 9.2: SKIP: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 9.2: SKIP: COMMA_K287_RXED_PLCWD",  "10",                      COMMA_K287_RXED_PLCWD,  test_failed);

  -- Test 9.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_SKIP_WORD & C_SKIP_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 9.3: SKIP: DATA_RX_PLCWD",          x"00000000" & x"00000000", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 9.3: SKIP: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 9.3: SKIP: DATA_RDY_PLCWD",         "00",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 9.3: SKIP: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 9.3: SKIP: COMMA_K287_RXED_PLCWD",  "11",                      COMMA_K287_RXED_PLCWD,  test_failed);

  --------------------------------------
  -- TEST 10: IDLE detect             --
  --------------------------------------
  -- Test 10.1: First word only
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678"& C_SKIP_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 10.1: IDLE: DATA_RX_PLCWD",          x"12345678"& x"00000000", DATA_RX_PLCWD,           test_failed);
  check_equal("Test 10.1: IDLE: VALID_K_CHARAC_PLCWD",   x"00",                    VALID_K_CHARAC_PLCWD,    test_failed);
  check_equal("Test 10.1: IDLE: DATA_RDY_PLCWD",         "10",                     DATA_RDY_PLCWD,          test_failed);
  check_equal("Test 10.1: IDLE: RX_NEW_WORD_PLCWD",      "11",                     RX_NEW_WORD_PLCWD,       test_failed);
  check_equal("Test 10.1: IDLE: COMMA_K287_RXED_PLCWD",  "01",                     COMMA_K287_RXED_PLCWD,   test_failed);

  -- Test 10.2: Second word only
  --------------------------------------
  DATA_RX_PLPL       <= C_IDLE_WORD & x"12345678";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 10.2: IDLE: DATA_RX_PLCWD",          x"00000000" & x"12345678", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 10.2: IDLE: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 10.2: IDLE: DATA_RDY_PLCWD",         "01",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 10.2: IDLE: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 10.2: IDLE: COMMA_K287_RXED_PLCWD",  "10",                      COMMA_K287_RXED_PLCWD,  test_failed);

  -- Test 10.3: 2 words
  --------------------------------------
  DATA_RX_PLPL       <= C_IDLE_WORD & C_IDLE_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 10.3: IDLE: DATA_RX_PLCWD",          x"00000000" & x"00000000", DATA_RX_PLCWD,          test_failed);
  check_equal("Test 10.3: IDLE: VALID_K_CHARAC_PLCWD",   x"00",                     VALID_K_CHARAC_PLCWD,   test_failed);
  check_equal("Test 10.3: IDLE: DATA_RDY_PLCWD",         "00",                      DATA_RDY_PLCWD,         test_failed);
  check_equal("Test 10.3: IDLE: RX_NEW_WORD_PLCWD",      "11",                      RX_NEW_WORD_PLCWD,      test_failed);
  check_equal("Test 10.3: IDLE: COMMA_K287_RXED_PLCWD",  "11",                      COMMA_K287_RXED_PLCWD,  test_failed);

  --------------------------------------
  -- TEST 11: ELSE                    --
  --------------------------------------
  ENABLE_TRANSM_DATA_PLIF <= '0';
  wait for 1 us;
  -- Test 11.1: 2 data words
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678" & x"9abcdef0";
  VALID_K_CHARAC_PLPL <= x"0" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 11.1: ELSE : DATA_RX_PLCWD",             x"00000000" & x"00000000", DATA_RX_PLCWD,             test_failed);
  check_equal("Test 11.1: ELSE : VALID_K_CHARAC_PLCWD",      x"00",                     VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 11.1: ELSE : DATA_RDY_PLCWD",            "00",                      DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 11.1: ELSE : RX_NEW_WORD_PLCWD",         "11",                      RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 11.1: ELSE : DETECTED_RXERR_WORD_PLCWD", "00",                      DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 11.2: First word only RXERR
  --------------------------------------
  DATA_RX_PLPL       <= x"12345678" & C_RXERR_WORD;
  VALID_K_CHARAC_PLPL <= x"0" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 11.2: ELSE : DATA_RX_PLCWD",             x"00000000" & x"00000000",  DATA_RX_PLCWD,             test_failed);
  check_equal("Test 11.2: ELSE : VALID_K_CHARAC_PLCWD",      x"00",                      VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 11.2: ELSE : DATA_RDY_PLCWD",            "00",                       DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 11.2: ELSE : RX_NEW_WORD_PLCWD",         "11",                       RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 11.2: ELSE : DETECTED_RXERR_WORD_PLCWD", "01",                       DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 11.3: Second word only RXERR
  --------------------------------------
  DATA_RX_PLPL       <= C_RXERR_WORD & x"9abcdef0";
  VALID_K_CHARAC_PLPL <= x"1" & x"0";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 11.3: ELSE : DATA_RX_PLCWD",             x"00000000" & x"00000000",  DATA_RX_PLCWD,             test_failed);
  check_equal("Test 11.3: ELSE : VALID_K_CHARAC_PLCWD",      x"00",                      VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 11.3: ELSE : DATA_RDY_PLCWD",            "00",                       DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 11.3: ELSE : RX_NEW_WORD_PLCWD",         "11",                       RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 11.1: ELSE : DETECTED_RXERR_WORD_PLCWD", "10",                       DETECTED_RXERR_WORD_PLCWD, test_failed);

  -- Test 11.4: 2 words RXERR
  --------------------------------------
  DATA_RX_PLPL       <= C_RXERR_WORD & C_RXERR_WORD;
  VALID_K_CHARAC_PLPL <= x"1" & x"1";
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check_equal("Test 11.4: ELSE : DATA_RX_PLCWD",             x"00000000" & x"00000000",   DATA_RX_PLCWD,             test_failed);
  check_equal("Test 11.4: ELSE : VALID_K_CHARAC_PLCWD",      x"00",                       VALID_K_CHARAC_PLCWD,      test_failed);
  check_equal("Test 11.4: ELSE : DATA_RDY_PLCWD",            "00",                        DATA_RDY_PLCWD,            test_failed);
  check_equal("Test 11.4: ELSE : RX_NEW_WORD_PLCWD",         "11",                        RX_NEW_WORD_PLCWD,         test_failed);
  check_equal("Test 11.4: ELSE : DETECTED_RXERR_WORD_PLCWD", "11",                        DETECTED_RXERR_WORD_PLCWD, test_failed);

  --------------------------------------
  -- TEST 12: NO SIGNAL detection     --
  --------------------------------------
  NO_SIGNAL_DETECTION_ENABLED_PLIF <= '1';
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check("Test 12: NO SIGNAL : NO_SIGNAL_PLCWD", '1', NO_SIGNAL_PLCWD, test_failed);

  NO_SIGNAL_DETECTION_ENABLED_PLIF <= '0';
  wait until falling_edge(CLK);
  wait until falling_edge(CLK);
  check("Test 12: NO SIGNAL : NO_SIGNAL_PLCWD", '0', NO_SIGNAL_PLCWD, test_failed);
  ------------------------------------------------------------
  --                       END TEST                         --
  ------------------------------------------------------------
  log_test_result(test_failed);

  wait;
end process;

end tb;