library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.data_link_lib.all;

entity data_link is
  generic(
    G_VC_NUM           : integer := 8                                                  --! Number of virtual channel
    );
  port(
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- Network layer AXI-Stream TX interface
    AXIS_ACLK_TX_DL        : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_TX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_TX_DL       : in  vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_TX_DL       : in  vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_TX_DL       : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_TX_DL      : in  std_logic_vector(G_VC_NUM downto 0);
    -- Network layer RX interface
    AXIS_ACLK_RX_DL        : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_RX_DL      : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_RX_DL       : out vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_RX_DL       : out vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_RX_DL       : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_RX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    -- Lane layer TX interface
    DATA_TX_PPL            : out  std_logic_vector(31 downto 00);     --! Data parallel to be send from Data-Link Layer
    CAPABILITY_TX_PPL      : out  std_logic_vector(07 downto 00);     --! Capability send on TX link in INIT3 control word
    NEW_DATA_TX_PPL        : out  std_logic;                          --! Flag to write data in FIFO TX
    VALID_K_CHARAC_TX_PPL  : out  std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TX_PPL vector
    FIFO_TX_FULL_PPL       : in   std_logic;                          --! Flag full of the FIFO TX
    -- Lane layer RX interface
    FIFO_RX_RD_EN_PPL      : out  std_logic;                          --! Flag to read data in FIFO RX
    DATA_RX_PPL            : in   std_logic_vector(31 downto 00);     --! Data parallel to be received to Data-Link Layer
    FIFO_RX_EMPTY_PPL      : in   std_logic;                          --! Flag EMPTY of the FIFO RX
    FIFO_RX_DATA_VALID_PPL : in   std_logic;                          --! Flag DATA_VALID of the FIFO RX
    VALID_K_CHARAC_RX_PPL  : in   std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TR_PPL vector
    FAR_END_CAPA_DL        : in   std_logic_vector(07 downto 00)     --! Capability field receive in INIT3 control word
    -- MIB  parameters interface
    INTERFACE_RESET_DL     : in std_logic;                            --! Reset the link and all configuration register of the Data Link layer
    LINK_RESET_DL          : in std_logic;                            --! Reset the link
    NACK_RST_EN_DL         : in std_logic;                            --! Enable automatic link reset on NACK reception
    NACK_RST_MODE_DL       : in std_logic;                            --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
    PAUSE_VC_DL            : in std_logic_vector(G_VC_NUM downto 0);         --! Pause the corresponding virtual channel after the end of current transmission
    CONTINUOUS_VC_DL       : in std_logic_vector(G_VC_NUM-1 downto 0);         --! Enable the corresponding virtual channel continuous mode   
    -- MIB  status interface
    SEQ_NUMBER_TX_DL        : out std_logic_vector(G_VC_NUM-1 downto 0);       --! SEQ_NUMBER in transmission
    SEQ_NUMBER_RX_DL        : out std_logic_vector(G_VC_NUM-1 downto 0);       --! SEQ_NUMBER in reception
    CREDIT_VC_DL            : out std_logic_vector(G_VC_NUM-1 downto 0);       --! Indicates if each corresponding far-end input buffer has credit
    FCT_CREDIT_OVERFLOW_DL  : out std_logic_vector(G_VC_NUM-1 downto 0);       --! Indicates overflow of each corresponding input buffer
    CRC_LONG_ERROR_DL       : out std_logic;                          --! CRC long error
    CRC_SHORT_ERROR_DL      : out std_logic;                          --! CRC short error
    FRAME_ERROR_DL          : out std_logic;                          --! Frame error
    SEQUENCE_ERROR_DL       : out std_logic;                          --! Sequence error
    FAR_END_LINK_RESET_DL   : out std_logic;                          --! Far-end link reset status
    FRAME_FINISHED_DL       : out std_logic_vector(G_VC_NUM downto 0);       --! Indicates that corresponding channel finished emitting a frame
    FRAME_TX_DL             : out std_logic_vector(G_VC_NUM downto 0);       --! Indicates that corresponding channel is emitting a frame
    DATA_COUNTER_TX_DL      : out std_logic_vector(6 downto 0);       --! Indicate the number of data transmitted in last frame emitted
    DATA_COUNTER_RX_DL      : out std_logic_vector(6 downto 0);       --! Indicate the number of data received in last frame received
    ACK_COUNTER_TX_DL       : out  std_logic_vector(2 downto 0);      --! ACK counter TX
    NACK_COUNTER_TX_DL      : out  std_logic_vector(2 downto 0);      --! NACK counter TX
    FCT_COUNTER_TX_DL       : out  std_logic_vector(3 downto 0);      --! FCT counter TX
    ACK_COUNTER_RX_DL       : out  std_logic_vector(2 downto 0);      --! ACK counter RX
    NACK_COUNTER_RX_DL      : out  std_logic_vector(2 downto 0);      --! NACK counter RX
    FCT_COUNTER_RX_DL       : out  std_logic_vector(3 downto 0);      --! FCT counter RX
    FULL_COUNTER_RX_DL      : out  std_logic_vector(1 downto 0);      --! FULL counter RX
    RETRY_COUNTER_RX_DL     : out  std_logic_vector(1 downto 0);      --! RETRY counter RX
    CURRENT_TIME_SLOT_DL    : out  std_logic_vector(7 downto 0)       --! Current time slot
  );
end data_link;

architecture Behavioral of data_link is
  -- Déclaration des composants
  component data_out_buff is
    port (
      RST_N                 : in  std_logic;                                    --! global reset
      CLK                   : in  std_logic;                                    --! Clock generated by GTY IP
      -- Link Reset
      LINK_RESET            : in std_logic;
      -- AXI-Stream interface
      S_AXIS_ACLK	          : in std_logic;
      S_AXIS_TREADY        	: out std_logic;
      S_AXIS_TDATA         	: in std_logic_vector(C_DATA_LENGTH-1 downto 0);
      S_AXIS_TUSER         	: in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      S_AXIS_TLAST         	: in std_logic;
      S_AXIS_TVALID        	: in std_logic;
      -- DOBUF interface
      VC_READY_DOBUF        : out  std_logic;
      DATA_DOBUF            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DOBUF  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      DATA_VALID_DOBUF      : out  std_logic;
      END_PACKET_DOBUF      : out  std_logic;
      VC_RD_EN_DMAC         : in   std_logic;
      --DDES interface
      M_VAL_DDES            : in std_logic_vector(C_M_SIZE-1 downto 0);
      FCT_FAR_END_DDES      : in std_logic;
      -- PPL interface
      LANE_ACTIVE_ST_PPL    : in std_logic;
      --MIB Interface
      FCT_CC_OVF_DOBUF      : out std_logic;
      VC_CONT_MODE_MIB      : in std_logic
    );
  end component;
  
  component data_mac is
    generic(
      G_VC_NUM           : integer := 8                                                  --! Number of virtual channel
      );
    port (
      RST_N              : in  std_logic;                                    --! global reset
      CLK                : in  std_logic;                                    --! Clock generated by GTY IP
      -- DERRM interface
      REQ_ACK_DERRM       : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      REQ_NACK_DERRM      : in  std_logic;
      TRANS_POL_FLG_DERRM : in  std_logic;
      REQ_ACK_DONE_DMAC   : out std_logic;
      -- DIBUF interface
      REQ_FCT_DIBUF       : in  std_logic_vector(G_VC_NUM-1 downto 0);                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      REQ_FCT_DONE_DIBUF  : out std_logic_vector(G_VC_NUM-1 downto 0);   
      -- DOBUF interface
      VC_READY_DOBUF      : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_DATA_DOBUF       : in  vc_data_array(G_VC_NUM-1 downto 0);
      VC_DATA_VALID_DOBUF : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_END_PACKET_DOBUF : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_RD_EN_DMAC       : out  std_logic_vector(G_VC_NUM-1 downto 0);
      -- MIB interface
      VC_PAUSE_MIB        : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_END_EMISSION_MIB : out std_logic_vector(G_VC_NUM-1 downto 0);
      VC_RUN_EMISSION_MIB : out std_logic_vector(G_VC_NUM-1 downto 0);
      -- DENC interface
      DATA_DMAC            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);  
      NEW_WORD_DMAC        : out std_logic;                                   
      NEW_PACKET_DMAC      : out std_logic;                                   
      END_PACKET_DMAC      : out std_logic;                                   
      TYPE_FRAME_DMAC      : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0); 
      VIRTUAL_CHANNEL_DMAC : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_TYPE_DMAC         : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_CHANNEL_DMAC      : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_STATUS_DMAC       : out std_logic_vector(2-1 downto 0);
      MULT_CHANNEL_DMAC    : out std_logic_vector(G_VC_NUM-1 downto 0);
      TRANS_POL_FLG_DMAC   : out std_logic;
      READY_DENC           : in std_logic
    );
  end component;
  component data_encpasulation IS
    generic (
        G_VC_NUM                       : INTEGER := 8                                                  --! Number of virtual channel
    );
    port (
      RST_N                            : IN  std_logic;                                    --! global reset
      CLK                              : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DMAC interface
      DATA_DMAC                        : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      NEW_WORD_DMAC                    : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      NEW_PACKET_DMAC                  : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      END_PACKET_DMAC                  : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      TYPE_FRAME_DMAC                  : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);                 --! Flag EMPTY of the FIFO RX
      VIRTUAL_CHANNEL_DMAC             : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_TYPE_DMAC                     : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_CHANNEL_DMAC                  : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_STATUS_DMAC                    : in std_logic_vector (2-1 downto 0);
      MULT_CHANNEL_DMAC                : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      -- DSCOM interface
      NEW_WORD_DENC                    : OUT  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DENC                        : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DENC              : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DENC                  : OUT  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);                 --! Flag EMPTY of the FIFO RX
      END_FRAME_DENC                   : OUT  std_logic
    );
  end component;

  component data_seq_compute IS
    port (
      RST_N                 : IN  std_logic;                                    --! global reset
      CLK                   : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DENC interface
      NEW_WORD_DENC         : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DENC        : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DENC   : IN  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DENC       : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DENC        : IN  std_logic;
      -- DCCOM interface
      NEW_WORD_DSCOM        : OUT  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DSCOM       : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DSCOM  : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DSCOM      : OUT  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DSCOM       : OUT  std_logic
    );
  end component;

  component data_crc_compute IS
    port (
      RST_N                 : IN  std_logic;                                    --! global reset
      CLK                   : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DSCOM interface
      NEW_WORD_DSCOM        : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DSCOM            : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DSCOM  : IN  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DSCOM      : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DSCOM       : IN  std_logic;
      -- FIFO_TX_LANE interface
      FIFO_FULL_TX_LANE     : IN  std_logic;
      VALID_K_CHARAC_DCCOM  : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      DATA_DCCOM            : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);    -- Data write bus
      NEW_WORD_DCCOM        : OUT  std_logic                                -- Write command
    );
  end component;
  signal LANE_ACTIVE_ST_PPL    : std_logic;
  -- DDES interface signals
  signal M_VAL_DDES            : vc_mult_array(G_VC_NUM-1 downto 0);
  signal FCT_FAR_END_DDES      : std_logic_vector(G_VC_NUM-1 downto 0);
  -- DOBUF interface signals
  signal VC_READY_DOBUF        : std_logic_vector(G_VC_NUM-1 downto 0);
  signal DATA_DOBUF            : vc_data_array(G_VC_NUM-1 downto 0);
  signal VALID_K_CHARAC_DOBUF  : vc_k_array(G_VC_NUM-1 downto 0);
  signal DATA_VALID_DOBUF      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal END_PACKET_DOBUF      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal FCT_CC_OVF_DOBUF      : std_logic_vector(G_VC_NUM-1 downto 0);
  
  -- DMAC interface signals
  signal DATA_DMAC                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal NEW_WORD_DMAC             : std_logic;
  signal NEW_PACKET_DMAC           : std_logic;
  signal END_PACKET_DMAC           : std_logic;
  signal TYPE_FRAME_DMAC           : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal VIRTUAL_CHANNEL_DMAC      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal BC_TYPE_DMAC              : std_logic_vector(G_VC_NUM-1 downto 0);
  signal BC_CHANNEL_DMAC           : std_logic_vector(G_VC_NUM-1 downto 0);
  signal BC_STATUS_DMAC            : std_logic_vector(2-1 downto 0);
  signal MULT_CHANNEL_DMAC         : std_logic_vector(G_VC_NUM-1 downto 0);
  signal REQ_ACK_DERRM             : std_logic;
  signal REQ_NACK_DERRM            : std_logic;
  signal TRANS_POL_FLG_DERRM       : std_logic;
  signal REQ_ACK_DONE_DMAC         : std_logic;
  signal REQ_FCT_DIBUF             : std_logic_vector(G_VC_NUM-1 downto 0);
  signal REQ_FCT_DONE_DIBUF        : std_logic_vector(G_VC_NUM-1 downto 0);   
  signal VC_RD_EN_DMAC             : std_logic_vector(G_VC_NUM-1 downto 0);
  signal VC_PAUSE_MIB              : std_logic_vector(G_VC_NUM-1 downto 0);
  signal VC_END_EMISSION_MIB       : std_logic_vector(G_VC_NUM-1 downto 0);
  signal VC_RUN_EMISSION_MIB       : std_logic_vector(G_VC_NUM-1 downto 0);

  -- DENC interface signals
  signal NEW_WORD_DENC             : std_logic;
  signal DATA_DENC                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal VALID_K_CHARAC_DENC       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal TYPE_FRAME_DENC           : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal END_FRAME_DENC            : std_logic;

  -- DSCOM interface signals
  signal NEW_WORD_DSCOM            : std_logic;
  signal DATA_DSCOM           : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal VALID_K_CHARAC_DSCOM      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal TYPE_FRAME_DSCOM          : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal END_FRAME_DSCOM           : std_logic;

  -- FIFO_TX_LANE interface signals
  signal FIFO_FULL_TX_LANE         : std_logic:='0';
  signal VALID_K_CHARAC_DCCOM      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal DATA_DCCOM                : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal NEW_WORD_DCCOM            : std_logic;

  -- DWI interface signals
  signal DATA_DWI                  : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal NEW_WORD_DWI              : std_logic;
  signal END_FRAME_DWI              : std_logic;
  signal SEQ_NUM_DWI                : std_logic_vector(7 downto 0);
  signal CRC_16B_DWI               : std_logic_vector(15 downto 0);
  signal CRC_8B_DWI                : std_logic_vector(7 downto 0);
  signal TYPE_FRAME_DWI            : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);

  -- CRC Check signals
  signal NEW_WORD_DCCHECK          : std_logic;
  signal DATA_DCCHECK         : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal SEQ_NUM_DCCHECK           : std_logic_vector(7 downto 0);
  signal END_FRAME_DCCHECK            : std_logic;
  signal CRC_ERR                   : std_logic;

  -- Sequence Check signals
  signal REC_POLARITY_FLG          : std_logic;
  signal TYPE_FRAME_DCCHECK        : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal SEQ_NUM_ERR               : std_logic;
  signal DATA_DSCHECK         : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal END_FRAME_DSCHECK               : std_logic;
  signal NEW_WORD_DSCHECK          : std_logic;
  signal FIFO_FULL                 : std_logic:='0';

  -- PHY PLUS LANE layer interface signals
  signal LINK_RESET                : std_logic;
  signal FRAME_ERR                 : std_logic;
  signal SEQ_ERR                    : std_logic;
  --MIB 
  signal VC_CONT_MODE_MIB         : std_logic_vector(G_VC_NUM-1 downto 0);

begin
    gen_data_out_buff: for i in 0 to G_VC_NUM-1 generate
      inst_data_out_buff: entity work.data_out_buff
          port map (
              RST_N                 => RST_N,
              CLK                   => CLK,
              LINK_RESET            => LINK_RESET,
              S_AXIS_ACLK           => AXIS_ACLK_TX_DL(i),
              S_AXIS_TREADY         => AXIS_TREADY_TX_DL(i),
              S_AXIS_TDATA          => AXIS_TDATA_TX_DL(i),
              S_AXIS_TUSER          => AXIS_TUSER_TX_DL(i),
              S_AXIS_TLAST          => AXIS_TLAST_TX_DL(i),
              S_AXIS_TVALID         => AXIS_TVALID_TX_DL(i),
              VC_READY_DOBUF        => VC_READY_DOBUF(i),
              DATA_DOBUF            => DATA_DOBUF(i),
              VALID_K_CHARAC_DOBUF  => VALID_K_CHARAC_DOBUF(i),
              DATA_VALID_DOBUF      => DATA_VALID_DOBUF(i),
              END_PACKET_DOBUF      => END_PACKET_DOBUF(i),
              VC_RD_EN_DMAC         => VC_RD_EN_DMAC(i),
              M_VAL_DDES            => M_VAL_DDES(i),
              FCT_FAR_END_DDES      => FCT_FAR_END_DDES(i),
              LANE_ACTIVE_ST_PPL    => LANE_ACTIVE_ST_PPL,
              FCT_CC_OVF_DOBUF      => FCT_CC_OVF_DOBUF(i),
              VC_CONT_MODE_MIB      => VC_CONT_MODE_MIB(i)
          );
  end generate;

  inst_data_mac: entity work.data_mac
    generic map (
        G_VC_NUM => G_VC_NUM
    );
    port map (
        RST_N                => RST_N,
        CLK                  => CLK,
        REQ_ACK_DERRM        => REQ_ACK_DERRM,
        REQ_NACK_DERRM       => REQ_NACK_DERRM,
        TRANS_POL_FLG_DERRM  => TRANS_POL_FLG_DERRM,
        REQ_ACK_DONE_DMAC    => REQ_ACK_DONE_DMAC,
        REQ_FCT_DIBUF        => REQ_FCT_DIBUF,
        VC_READY_DOBUF       => VC_READY_DOBUF,
        VC_DATA_DOBUF        => VC_DATA_DOBUF,
        VC_DATA_VALID_DOBUF  => VC_DATA_VALID_DOBUF,
        VC_RD_EN_DMAC        => VC_RD_EN_DMAC,
        VC_PAUSE_MIB         => VC_PAUSE_MIB,
        VC_END_EMISSION_MIB  => VC_END_EMISSION_MIB,
        VC_END_PACKET_DOBUF  => VC_END_PACKET_DOBUF,
        VC_RUN_EMISSION_MIB  => VC_RUN_EMISSION_MIB,
        DATA_DMAC            => DATA_DMAC,
        NEW_WORD_DMAC        => NEW_WORD_DMAC,
        NEW_PACKET_DMAC      => NEW_PACKET_DMAC,
        END_PACKET_DMAC      => END_PACKET_DMAC,
        TYPE_FRAME_DMAC      => TYPE_FRAME_DMAC,
        VIRTUAL_CHANNEL_DMAC => VIRTUAL_CHANNEL_DMAC,
        BC_TYPE_DMAC         => BC_TYPE_DMAC,
        BC_CHANNEL_DMAC      => BC_CHANNEL_DMAC,
        BC_STATUS_DMAC       => BC_STATUS_DMAC,
        MULT_CHANNEL_DMAC    => MULT_CHANNEL_DMAC,
        TRANS_POL_FLG_DMAC   => TRANS_POL_FLG_DMAC,
        READY_DENC           => READY_DENC
    );
  
  inst_data_encpasulation: entity work.data_encpasulation
      generic map (
          G_VC_NUM => G_VC_NUM
      );
      port map (
          RST_N                 => RST_N,
          CLK                   => CLK,
          DATA_DMAC             => DATA_DMAC,
          NEW_WORD_DMAC         => NEW_WORD_DMAC,
          NEW_PACKET_DMAC       => NEW_PACKET_DMAC,
          END_PACKET_DMAC       => END_PACKET_DMAC,
          TYPE_FRAME_DMAC       => TYPE_FRAME_DMAC,
          VIRTUAL_CHANNEL_DMAC  => VIRTUAL_CHANNEL_DMAC,
          BC_TYPE_DMAC          => BC_TYPE_DMAC,
          BC_CHANNEL_DMAC       => BC_CHANNEL_DMAC,
          BC_STATUS_DMAC        => BC_STATUS_DMAC,
          MULT_CHANNEL_DMAC     => MULT_CHANNEL_DMAC,
          NEW_WORD_DENC         => NEW_WORD_DENC,
          DATA_DENC             => DATA_DENC,
          VALID_K_CHARAC_DENC   => VALID_K_CHARAC_DENC,
          TYPE_FRAME_DENC       => TYPE_FRAME_DENC,
          END_FRAME_DENC        => END_FRAME_DENC
      );

    inst_data_seq_compute: entity work.data_seq_compute
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            NEW_WORD_DENC         => NEW_WORD_DENC,
            DATA_DENC        => DATA_DENC,
            VALID_K_CHARAC_DENC   => VALID_K_CHARAC_DENC,
            TYPE_FRAME_DENC       => TYPE_FRAME_DENC,
            END_FRAME_DENC        => END_FRAME_DENC,
            NEW_WORD_DSCOM        => NEW_WORD_DSCOM,
            DATA_DSCOM       => DATA_DSCOM,
            VALID_K_CHARAC_DSCOM  => VALID_K_CHARAC_DSCOM,
            TYPE_FRAME_DSCOM      => TYPE_FRAME_DSCOM,
            END_FRAME_DSCOM       => END_FRAME_DSCOM
        );

    inst_data_crc_compute: entity work.data_crc_compute
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            NEW_WORD_DSCOM        => NEW_WORD_DSCOM,
            DATA_DSCOM            => DATA_DSCOM,
            VALID_K_CHARAC_DSCOM  => VALID_K_CHARAC_DSCOM,
            TYPE_FRAME_DSCOM      => TYPE_FRAME_DSCOM,
            END_FRAME_DSCOM       => END_FRAME_DSCOM,
            FIFO_FULL_TX_LANE     => FIFO_FULL_TX_LANE,
            VALID_K_CHARAC_DCCOM  => VALID_K_CHARAC_DCCOM,
            DATA_DCCOM            => DATA_DCCOM,
            NEW_WORD_DCCOM        => NEW_WORD_DCCOM
        );

end Behavioral;
