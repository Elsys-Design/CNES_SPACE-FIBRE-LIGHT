// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_X5PHIO_XCVR_X2_DEFINES_VH
`else
`define B_X5PHIO_XCVR_X2_DEFINES_VH

// Look-up table parameters
//

`define X5PHIO_XCVR_X2_ADDR_N  156
`define X5PHIO_XCVR_X2_ADDR_SZ 32
`define X5PHIO_XCVR_X2_DATA_SZ 152

// Attribute addresses
//

`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_POL_M    32'h00000000
`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_POL_S    32'h00000001
`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_VALUE_M    32'h00000002
`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_VALUE_M_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_VALUE_S    32'h00000003
`define X5PHIO_XCVR_X2__ADL_H1ME_OFST_VALUE_S_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_POL_M    32'h00000004
`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_POL_S    32'h00000005
`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_VALUE_M    32'h00000006
`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_VALUE_M_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_VALUE_S    32'h00000007
`define X5PHIO_XCVR_X2__ADL_H1MO_OFST_VALUE_S_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_POL_M    32'h00000008
`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_POL_S    32'h00000009
`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_VALUE_M    32'h0000000a
`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_VALUE_M_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_VALUE_S    32'h0000000b
`define X5PHIO_XCVR_X2__ADL_H1PE_OFST_VALUE_S_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_POL_M    32'h0000000c
`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_POL_S    32'h0000000d
`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_VALUE_M    32'h0000000e
`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_VALUE_M_SZ 4

`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_VALUE_S    32'h0000000f
`define X5PHIO_XCVR_X2__ADL_H1PO_OFST_VALUE_S_SZ 4

`define X5PHIO_XCVR_X2__APBCLK_FREQ    32'h00000010
`define X5PHIO_XCVR_X2__APBCLK_FREQ_SZ 9

`define X5PHIO_XCVR_X2__CASCADE_IDL_M    32'h00000011
`define X5PHIO_XCVR_X2__CASCADE_IDL_M_SZ 96

`define X5PHIO_XCVR_X2__CASCADE_IDL_S    32'h00000012
`define X5PHIO_XCVR_X2__CASCADE_IDL_S_SZ 96

`define X5PHIO_XCVR_X2__CASCADE_ODL_M    32'h00000013
`define X5PHIO_XCVR_X2__CASCADE_ODL_M_SZ 104

`define X5PHIO_XCVR_X2__CASCADE_ODL_S    32'h00000014
`define X5PHIO_XCVR_X2__CASCADE_ODL_S_SZ 104

`define X5PHIO_XCVR_X2__CCIO_EN_M    32'h00000015
`define X5PHIO_XCVR_X2__CCIO_EN_M_SZ 40

`define X5PHIO_XCVR_X2__CCIO_EN_S    32'h00000016
`define X5PHIO_XCVR_X2__CCIO_EN_S_SZ 40

`define X5PHIO_XCVR_X2__CLOCK_FREQ    32'h00000017
`define X5PHIO_XCVR_X2__CLOCK_FREQ_SZ 13

`define X5PHIO_XCVR_X2__CONTINUOUS_DQS    32'h00000018
`define X5PHIO_XCVR_X2__CONTINUOUS_DQS_SZ 40

`define X5PHIO_XCVR_X2__CPHY_MODE_CTRL    32'h00000019
`define X5PHIO_XCVR_X2__CPHY_MODE_CTRL_SZ 1

`define X5PHIO_XCVR_X2__CPHY_TERM_M    32'h0000001a
`define X5PHIO_XCVR_X2__CPHY_TERM_M_SZ 40

`define X5PHIO_XCVR_X2__CPHY_TERM_S    32'h0000001b
`define X5PHIO_XCVR_X2__CPHY_TERM_S_SZ 40

`define X5PHIO_XCVR_X2__CTLE_EQ_M    32'h0000001c
`define X5PHIO_XCVR_X2__CTLE_EQ_M_SZ 112

`define X5PHIO_XCVR_X2__CTLE_EQ_S    32'h0000001d
`define X5PHIO_XCVR_X2__CTLE_EQ_S_SZ 112

`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_POL_M    32'h0000001e
`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_POL_S    32'h0000001f
`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_VAL_M    32'h00000020
`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_VAL_S    32'h00000021
`define X5PHIO_XCVR_X2__CTLE_H1M_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_POL_M    32'h00000022
`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_POL_S    32'h00000023
`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_VAL_M    32'h00000024
`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_VAL_S    32'h00000025
`define X5PHIO_XCVR_X2__CTLE_H1P_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__CTLE_OFST_M    32'h00000026
`define X5PHIO_XCVR_X2__CTLE_OFST_M_SZ 128

`define X5PHIO_XCVR_X2__CTLE_OFST_S    32'h00000027
`define X5PHIO_XCVR_X2__CTLE_OFST_S_SZ 128

`define X5PHIO_XCVR_X2__DFE_EQ_M    32'h00000028
`define X5PHIO_XCVR_X2__DFE_EQ_M_SZ 120

`define X5PHIO_XCVR_X2__DFE_EQ_S    32'h00000029
`define X5PHIO_XCVR_X2__DFE_EQ_S_SZ 120

`define X5PHIO_XCVR_X2__DFE_H2_NEG_POL_M    32'h0000002a
`define X5PHIO_XCVR_X2__DFE_H2_NEG_POL_M_SZ 1

`define X5PHIO_XCVR_X2__DFE_H2_NEG_POL_S    32'h0000002b
`define X5PHIO_XCVR_X2__DFE_H2_NEG_POL_S_SZ 1

`define X5PHIO_XCVR_X2__DFE_H2_TAP_WEIGHT_M    32'h0000002c
`define X5PHIO_XCVR_X2__DFE_H2_TAP_WEIGHT_M_SZ 5

`define X5PHIO_XCVR_X2__DFE_H2_TAP_WEIGHT_S    32'h0000002d
`define X5PHIO_XCVR_X2__DFE_H2_TAP_WEIGHT_S_SZ 5

`define X5PHIO_XCVR_X2__DFE_H3_NEG_POL_M    32'h0000002e
`define X5PHIO_XCVR_X2__DFE_H3_NEG_POL_M_SZ 1

`define X5PHIO_XCVR_X2__DFE_H3_NEG_POL_S    32'h0000002f
`define X5PHIO_XCVR_X2__DFE_H3_NEG_POL_S_SZ 1

`define X5PHIO_XCVR_X2__DFE_H3_TAP_WEIGHT_M    32'h00000030
`define X5PHIO_XCVR_X2__DFE_H3_TAP_WEIGHT_M_SZ 5

`define X5PHIO_XCVR_X2__DFE_H3_TAP_WEIGHT_S    32'h00000031
`define X5PHIO_XCVR_X2__DFE_H3_TAP_WEIGHT_S_SZ 5

`define X5PHIO_XCVR_X2__DFE_H4_NEG_POL_M    32'h00000032
`define X5PHIO_XCVR_X2__DFE_H4_NEG_POL_M_SZ 1

`define X5PHIO_XCVR_X2__DFE_H4_NEG_POL_S    32'h00000033
`define X5PHIO_XCVR_X2__DFE_H4_NEG_POL_S_SZ 1

`define X5PHIO_XCVR_X2__DFE_H4_TAP_WEIGHT_M    32'h00000034
`define X5PHIO_XCVR_X2__DFE_H4_TAP_WEIGHT_M_SZ 4

`define X5PHIO_XCVR_X2__DFE_H4_TAP_WEIGHT_S    32'h00000035
`define X5PHIO_XCVR_X2__DFE_H4_TAP_WEIGHT_S_SZ 4

`define X5PHIO_XCVR_X2__DFE_INIT_M    32'h00000036
`define X5PHIO_XCVR_X2__DFE_INIT_M_SZ 40

`define X5PHIO_XCVR_X2__DFE_INIT_S    32'h00000037
`define X5PHIO_XCVR_X2__DFE_INIT_S_SZ 40

`define X5PHIO_XCVR_X2__DIFF_PIN_SWAP    32'h00000038
`define X5PHIO_XCVR_X2__DIFF_PIN_SWAP_SZ 40

`define X5PHIO_XCVR_X2__DIFF_SLAVE_RX_EN    32'h00000039
`define X5PHIO_XCVR_X2__DIFF_SLAVE_RX_EN_SZ 40

`define X5PHIO_XCVR_X2__DIFF_TERM    32'h0000003a
`define X5PHIO_XCVR_X2__DIFF_TERM_SZ 40

`define X5PHIO_XCVR_X2__DIV64CLK_EN    32'h0000003b
`define X5PHIO_XCVR_X2__DIV64CLK_EN_SZ 40

`define X5PHIO_XCVR_X2__DQS_ANA_DETECTION_M    32'h0000003c
`define X5PHIO_XCVR_X2__DQS_ANA_DETECTION_M_SZ 40

`define X5PHIO_XCVR_X2__DQS_ANA_DETECTION_S    32'h0000003d
`define X5PHIO_XCVR_X2__DQS_ANA_DETECTION_S_SZ 40

`define X5PHIO_XCVR_X2__DQS_BIAS_M    32'h0000003e
`define X5PHIO_XCVR_X2__DQS_BIAS_M_SZ 40

`define X5PHIO_XCVR_X2__DQS_BIAS_S    32'h0000003f
`define X5PHIO_XCVR_X2__DQS_BIAS_S_SZ 40

`define X5PHIO_XCVR_X2__DRIVE_M    32'h00000040
`define X5PHIO_XCVR_X2__DRIVE_M_SZ 5

`define X5PHIO_XCVR_X2__DRIVE_S    32'h00000041
`define X5PHIO_XCVR_X2__DRIVE_S_SZ 5

`define X5PHIO_XCVR_X2__DYNAMIC_DCI_TS_0    32'h00000042
`define X5PHIO_XCVR_X2__DYNAMIC_DCI_TS_0_SZ 40

`define X5PHIO_XCVR_X2__DYNAMIC_DCI_TS_1    32'h00000043
`define X5PHIO_XCVR_X2__DYNAMIC_DCI_TS_1_SZ 40

`define X5PHIO_XCVR_X2__EN_OMUX    32'h00000044
`define X5PHIO_XCVR_X2__EN_OMUX_SZ 40

`define X5PHIO_XCVR_X2__IO_TYPE_M    32'h00000045
`define X5PHIO_XCVR_X2__IO_TYPE_M_SZ 80

`define X5PHIO_XCVR_X2__IO_TYPE_S    32'h00000046
`define X5PHIO_XCVR_X2__IO_TYPE_S_SZ 80

`define X5PHIO_XCVR_X2__ISTANDARD_M    32'h00000047
`define X5PHIO_XCVR_X2__ISTANDARD_M_SZ 48

`define X5PHIO_XCVR_X2__ISTANDARD_S    32'h00000048
`define X5PHIO_XCVR_X2__ISTANDARD_S_SZ 48

`define X5PHIO_XCVR_X2__LL_2TO1_MODE_0    32'h00000049
`define X5PHIO_XCVR_X2__LL_2TO1_MODE_0_SZ 40

`define X5PHIO_XCVR_X2__LL_2TO1_MODE_1    32'h0000004a
`define X5PHIO_XCVR_X2__LL_2TO1_MODE_1_SZ 40

`define X5PHIO_XCVR_X2__MIPI_ALPRX_EN_M    32'h0000004b
`define X5PHIO_XCVR_X2__MIPI_ALPRX_EN_M_SZ 40

`define X5PHIO_XCVR_X2__MIPI_ALPRX_EN_S    32'h0000004c
`define X5PHIO_XCVR_X2__MIPI_ALPRX_EN_S_SZ 40

`define X5PHIO_XCVR_X2__MIPI_ALPTX_EN_M    32'h0000004d
`define X5PHIO_XCVR_X2__MIPI_ALPTX_EN_M_SZ 40

`define X5PHIO_XCVR_X2__MIPI_ALPTX_EN_S    32'h0000004e
`define X5PHIO_XCVR_X2__MIPI_ALPTX_EN_S_SZ 40

`define X5PHIO_XCVR_X2__MIPI_CPHY_PAD_M    32'h0000004f
`define X5PHIO_XCVR_X2__MIPI_CPHY_PAD_M_SZ 120

`define X5PHIO_XCVR_X2__MIPI_CPHY_PAD_S    32'h00000050
`define X5PHIO_XCVR_X2__MIPI_CPHY_PAD_S_SZ 120

`define X5PHIO_XCVR_X2__ODLY_SRC_M    32'h00000051
`define X5PHIO_XCVR_X2__ODLY_SRC_M_SZ 2

`define X5PHIO_XCVR_X2__ODLY_SRC_S    32'h00000052
`define X5PHIO_XCVR_X2__ODLY_SRC_S_SZ 2

`define X5PHIO_XCVR_X2__OSTANDARD_M    32'h00000053
`define X5PHIO_XCVR_X2__OSTANDARD_M_SZ 48

`define X5PHIO_XCVR_X2__OSTANDARD_S    32'h00000054
`define X5PHIO_XCVR_X2__OSTANDARD_S_SZ 48

`define X5PHIO_XCVR_X2__PHY2IOB_T_0    32'h00000055
`define X5PHIO_XCVR_X2__PHY2IOB_T_0_SZ 40

`define X5PHIO_XCVR_X2__PHY2IOB_T_1    32'h00000056
`define X5PHIO_XCVR_X2__PHY2IOB_T_1_SZ 40

`define X5PHIO_XCVR_X2__PHY2XCV_LATENCY    32'h00000057
`define X5PHIO_XCVR_X2__PHY2XCV_LATENCY_SZ 4

`define X5PHIO_XCVR_X2__RD_CTL_MUXSEL    32'h00000058
`define X5PHIO_XCVR_X2__RD_CTL_MUXSEL_SZ 8

`define X5PHIO_XCVR_X2__RIUCLK_DBLR_BYPASS    32'h00000059
`define X5PHIO_XCVR_X2__RIUCLK_DBLR_BYPASS_SZ 40

`define X5PHIO_XCVR_X2__ROUTETHRU_0    32'h0000005a
`define X5PHIO_XCVR_X2__ROUTETHRU_0_SZ 40

`define X5PHIO_XCVR_X2__ROUTETHRU_1    32'h0000005b
`define X5PHIO_XCVR_X2__ROUTETHRU_1_SZ 40

`define X5PHIO_XCVR_X2__RX2TX_LOOPBACK_M    32'h0000005c
`define X5PHIO_XCVR_X2__RX2TX_LOOPBACK_M_SZ 40

`define X5PHIO_XCVR_X2__RX2TX_LOOPBACK_S    32'h0000005d
`define X5PHIO_XCVR_X2__RX2TX_LOOPBACK_S_SZ 40

`define X5PHIO_XCVR_X2__RX_CLOCK    32'h0000005e
`define X5PHIO_XCVR_X2__RX_CLOCK_SZ 88

`define X5PHIO_XCVR_X2__RX_CLOCK_ALIGN_M    32'h0000005f
`define X5PHIO_XCVR_X2__RX_CLOCK_ALIGN_M_SZ 152

`define X5PHIO_XCVR_X2__RX_CLOCK_ALIGN_S    32'h00000060
`define X5PHIO_XCVR_X2__RX_CLOCK_ALIGN_S_SZ 152

`define X5PHIO_XCVR_X2__RX_DATA_WIDTH_M    32'h00000061
`define X5PHIO_XCVR_X2__RX_DATA_WIDTH_M_SZ 5

`define X5PHIO_XCVR_X2__RX_DATA_WIDTH_S    32'h00000062
`define X5PHIO_XCVR_X2__RX_DATA_WIDTH_S_SZ 5

`define X5PHIO_XCVR_X2__RX_GATING    32'h00000063
`define X5PHIO_XCVR_X2__RX_GATING_SZ 56

`define X5PHIO_XCVR_X2__RX_LOAD_DLY    32'h00000064
`define X5PHIO_XCVR_X2__RX_LOAD_DLY_SZ 2

`define X5PHIO_XCVR_X2__SA_H1ME_OFST_POL_M    32'h00000065
`define X5PHIO_XCVR_X2__SA_H1ME_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__SA_H1ME_OFST_POL_S    32'h00000066
`define X5PHIO_XCVR_X2__SA_H1ME_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__SA_H1ME_OFST_VAL_M    32'h00000067
`define X5PHIO_XCVR_X2__SA_H1ME_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__SA_H1ME_OFST_VAL_S    32'h00000068
`define X5PHIO_XCVR_X2__SA_H1ME_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__SA_H1MO_OFST_POL_M    32'h00000069
`define X5PHIO_XCVR_X2__SA_H1MO_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__SA_H1MO_OFST_POL_S    32'h0000006a
`define X5PHIO_XCVR_X2__SA_H1MO_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__SA_H1MO_OFST_VAL_M    32'h0000006b
`define X5PHIO_XCVR_X2__SA_H1MO_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__SA_H1MO_OFST_VAL_S    32'h0000006c
`define X5PHIO_XCVR_X2__SA_H1MO_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__SA_H1PE_OFST_POL_M    32'h0000006d
`define X5PHIO_XCVR_X2__SA_H1PE_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__SA_H1PE_OFST_POL_S    32'h0000006e
`define X5PHIO_XCVR_X2__SA_H1PE_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__SA_H1PE_OFST_VAL_M    32'h0000006f
`define X5PHIO_XCVR_X2__SA_H1PE_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__SA_H1PE_OFST_VAL_S    32'h00000070
`define X5PHIO_XCVR_X2__SA_H1PE_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__SA_H1PO_OFST_POL_M    32'h00000071
`define X5PHIO_XCVR_X2__SA_H1PO_OFST_POL_M_SZ 1

`define X5PHIO_XCVR_X2__SA_H1PO_OFST_POL_S    32'h00000072
`define X5PHIO_XCVR_X2__SA_H1PO_OFST_POL_S_SZ 1

`define X5PHIO_XCVR_X2__SA_H1PO_OFST_VAL_M    32'h00000073
`define X5PHIO_XCVR_X2__SA_H1PO_OFST_VAL_M_SZ 6

`define X5PHIO_XCVR_X2__SA_H1PO_OFST_VAL_S    32'h00000074
`define X5PHIO_XCVR_X2__SA_H1PO_OFST_VAL_S_SZ 6

`define X5PHIO_XCVR_X2__SA_OFST_CAL_M    32'h00000075
`define X5PHIO_XCVR_X2__SA_OFST_CAL_M_SZ 112

`define X5PHIO_XCVR_X2__SA_OFST_CAL_S    32'h00000076
`define X5PHIO_XCVR_X2__SA_OFST_CAL_S_SZ 112

`define X5PHIO_XCVR_X2__SIM_VERSION    32'h00000077
`define X5PHIO_XCVR_X2__SIM_VERSION_SZ 2

`define X5PHIO_XCVR_X2__SLEW_M    32'h00000078
`define X5PHIO_XCVR_X2__SLEW_M_SZ 48

`define X5PHIO_XCVR_X2__SLEW_S    32'h00000079
`define X5PHIO_XCVR_X2__SLEW_S_SZ 48

`define X5PHIO_XCVR_X2__SLV_WRLVL_MODE    32'h0000007a
`define X5PHIO_XCVR_X2__SLV_WRLVL_MODE_SZ 40

`define X5PHIO_XCVR_X2__TX0_ANALOG_SPARE0    32'h0000007b
`define X5PHIO_XCVR_X2__TX0_ANALOG_SPARE0_SZ 8

`define X5PHIO_XCVR_X2__TX0_DIG_SPARE0    32'h0000007c
`define X5PHIO_XCVR_X2__TX0_DIG_SPARE0_SZ 8

`define X5PHIO_XCVR_X2__TX0_ODLY_CASC_EN    32'h0000007d
`define X5PHIO_XCVR_X2__TX0_ODLY_CASC_EN_SZ 40

`define X5PHIO_XCVR_X2__TX0_OUTPUT_PHASE_90    32'h0000007e
`define X5PHIO_XCVR_X2__TX0_OUTPUT_PHASE_90_SZ 40

`define X5PHIO_XCVR_X2__TX1_ANALOG_SPARE0    32'h0000007f
`define X5PHIO_XCVR_X2__TX1_ANALOG_SPARE0_SZ 8

`define X5PHIO_XCVR_X2__TX1_DIG_SPARE0    32'h00000080
`define X5PHIO_XCVR_X2__TX1_DIG_SPARE0_SZ 8

`define X5PHIO_XCVR_X2__TX1_ODLY_CASC_EN    32'h00000081
`define X5PHIO_XCVR_X2__TX1_ODLY_CASC_EN_SZ 40

`define X5PHIO_XCVR_X2__TX1_OUTPUT_PHASE_90    32'h00000082
`define X5PHIO_XCVR_X2__TX1_OUTPUT_PHASE_90_SZ 40

`define X5PHIO_XCVR_X2__TX2RX_PREDRV_LOOPBACK_M    32'h00000083
`define X5PHIO_XCVR_X2__TX2RX_PREDRV_LOOPBACK_M_SZ 40

`define X5PHIO_XCVR_X2__TX2RX_PREDRV_LOOPBACK_S    32'h00000084
`define X5PHIO_XCVR_X2__TX2RX_PREDRV_LOOPBACK_S_SZ 40

`define X5PHIO_XCVR_X2__TX2RX_RETIMER_LOOPBACK_M    32'h00000085
`define X5PHIO_XCVR_X2__TX2RX_RETIMER_LOOPBACK_M_SZ 40

`define X5PHIO_XCVR_X2__TX2RX_RETIMER_LOOPBACK_S    32'h00000086
`define X5PHIO_XCVR_X2__TX2RX_RETIMER_LOOPBACK_S_SZ 40

`define X5PHIO_XCVR_X2__TX_DATA_WIDTH    32'h00000087
`define X5PHIO_XCVR_X2__TX_DATA_WIDTH_SZ 5

`define X5PHIO_XCVR_X2__TX_DRV_HP_EN_M    32'h00000088
`define X5PHIO_XCVR_X2__TX_DRV_HP_EN_M_SZ 40

`define X5PHIO_XCVR_X2__TX_DRV_HP_EN_S    32'h00000089
`define X5PHIO_XCVR_X2__TX_DRV_HP_EN_S_SZ 40

`define X5PHIO_XCVR_X2__TX_INIT_0    32'h0000008a
`define X5PHIO_XCVR_X2__TX_INIT_0_SZ 40

`define X5PHIO_XCVR_X2__TX_INIT_1    32'h0000008b
`define X5PHIO_XCVR_X2__TX_INIT_1_SZ 40

`define X5PHIO_XCVR_X2__TX_INIT_T    32'h0000008c
`define X5PHIO_XCVR_X2__TX_INIT_T_SZ 40

`define X5PHIO_XCVR_X2__USE_IBUFDISABLE_M    32'h0000008d
`define X5PHIO_XCVR_X2__USE_IBUFDISABLE_M_SZ 144

`define X5PHIO_XCVR_X2__USE_IBUFDISABLE_S    32'h0000008e
`define X5PHIO_XCVR_X2__USE_IBUFDISABLE_S_SZ 144

`define X5PHIO_XCVR_X2__VREF_H1M_PER_OCTAD_M    32'h0000008f
`define X5PHIO_XCVR_X2__VREF_H1M_PER_OCTAD_M_SZ 1

`define X5PHIO_XCVR_X2__VREF_H1M_PER_OCTAD_S    32'h00000090
`define X5PHIO_XCVR_X2__VREF_H1M_PER_OCTAD_S_SZ 1

`define X5PHIO_XCVR_X2__VREF_H1M_VALUE_M    32'h00000091
`define X5PHIO_XCVR_X2__VREF_H1M_VALUE_M_SZ 10

`define X5PHIO_XCVR_X2__VREF_H1M_VALUE_S    32'h00000092
`define X5PHIO_XCVR_X2__VREF_H1M_VALUE_S_SZ 10

`define X5PHIO_XCVR_X2__VREF_H1P_PER_OCTAD_M    32'h00000093
`define X5PHIO_XCVR_X2__VREF_H1P_PER_OCTAD_M_SZ 1

`define X5PHIO_XCVR_X2__VREF_H1P_PER_OCTAD_S    32'h00000094
`define X5PHIO_XCVR_X2__VREF_H1P_PER_OCTAD_S_SZ 1

`define X5PHIO_XCVR_X2__VREF_H1P_VALUE_M    32'h00000095
`define X5PHIO_XCVR_X2__VREF_H1P_VALUE_M_SZ 10

`define X5PHIO_XCVR_X2__VREF_H1P_VALUE_S    32'h00000096
`define X5PHIO_XCVR_X2__VREF_H1P_VALUE_S_SZ 10

`define X5PHIO_XCVR_X2__WR_CTL_MUXSEL    32'h00000097
`define X5PHIO_XCVR_X2__WR_CTL_MUXSEL_SZ 8

`define X5PHIO_XCVR_X2__WR_DQ0_MUXSEL    32'h00000098
`define X5PHIO_XCVR_X2__WR_DQ0_MUXSEL_SZ 8

`define X5PHIO_XCVR_X2__WR_DQ1_MUXSEL    32'h00000099
`define X5PHIO_XCVR_X2__WR_DQ1_MUXSEL_SZ 8

`define X5PHIO_XCVR_X2__WR_EN0_MUXSEL    32'h0000009a
`define X5PHIO_XCVR_X2__WR_EN0_MUXSEL_SZ 8

`define X5PHIO_XCVR_X2__WR_EN1_MUXSEL    32'h0000009b
`define X5PHIO_XCVR_X2__WR_EN1_MUXSEL_SZ 8

`endif  // B_X5PHIO_XCVR_X2_DEFINES_VH