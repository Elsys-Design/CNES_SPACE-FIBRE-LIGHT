`include "B_OSERDESE3_defines.vh"

reg [`OSERDESE3_DATA_SZ-1:0] ATTR [0:`OSERDESE3_ADDR_N-1];
reg [`OSERDESE3__DATA_WIDTH_SZ-1:0] DATA_WIDTH_REG = DATA_WIDTH;
reg INIT_REG = INIT;
reg IS_CLKDIV_INVERTED_REG = IS_CLKDIV_INVERTED;
reg IS_CLK_INVERTED_REG = IS_CLK_INVERTED;
reg IS_RST_INVERTED_REG = IS_RST_INVERTED;
reg [`OSERDESE3__ODDR_MODE_SZ:1] ODDR_MODE_REG = ODDR_MODE;
reg [`OSERDESE3__OSERDES_D_BYPASS_SZ:1] OSERDES_D_BYPASS_REG = OSERDES_D_BYPASS;
reg [`OSERDESE3__OSERDES_T_BYPASS_SZ:1] OSERDES_T_BYPASS_REG = OSERDES_T_BYPASS;
reg [`OSERDESE3__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
real SIM_VERSION_REG = SIM_VERSION;

initial begin
  ATTR[`OSERDESE3__DATA_WIDTH] = DATA_WIDTH;
  ATTR[`OSERDESE3__INIT] = INIT;
  ATTR[`OSERDESE3__IS_CLKDIV_INVERTED] = IS_CLKDIV_INVERTED;
  ATTR[`OSERDESE3__IS_CLK_INVERTED] = IS_CLK_INVERTED;
  ATTR[`OSERDESE3__IS_RST_INVERTED] = IS_RST_INVERTED;
  ATTR[`OSERDESE3__ODDR_MODE] = ODDR_MODE;
  ATTR[`OSERDESE3__OSERDES_D_BYPASS] = OSERDES_D_BYPASS;
  ATTR[`OSERDESE3__OSERDES_T_BYPASS] = OSERDES_T_BYPASS;
  ATTR[`OSERDESE3__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`OSERDESE3__SIM_VERSION] = $realtobits(SIM_VERSION);
end

always @(trig_attr) begin
  DATA_WIDTH_REG = ATTR[`OSERDESE3__DATA_WIDTH];
  INIT_REG = ATTR[`OSERDESE3__INIT];
  IS_CLKDIV_INVERTED_REG = ATTR[`OSERDESE3__IS_CLKDIV_INVERTED];
  IS_CLK_INVERTED_REG = ATTR[`OSERDESE3__IS_CLK_INVERTED];
  IS_RST_INVERTED_REG = ATTR[`OSERDESE3__IS_RST_INVERTED];
  ODDR_MODE_REG = ATTR[`OSERDESE3__ODDR_MODE];
  OSERDES_D_BYPASS_REG = ATTR[`OSERDESE3__OSERDES_D_BYPASS];
  OSERDES_T_BYPASS_REG = ATTR[`OSERDESE3__OSERDES_T_BYPASS];
  SIM_DEVICE_REG = ATTR[`OSERDESE3__SIM_DEVICE];
  SIM_VERSION_REG = $bitstoreal(ATTR[`OSERDESE3__SIM_VERSION]);
end

// procedures to override, read attribute values

task write_attr;
  input  [`OSERDESE3_ADDR_SZ-1:0] addr;
  input  [`OSERDESE3_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`OSERDESE3_DATA_SZ-1:0] read_attr;
  input  [`OSERDESE3_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
