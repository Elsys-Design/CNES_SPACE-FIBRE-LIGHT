// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC2_NMU128_DEFINES_VH
`else
`define B_NOC2_NMU128_DEFINES_VH

// Look-up table parameters
//

`define NOC2_NMU128_ADDR_N  295
`define NOC2_NMU128_ADDR_SZ 32
`define NOC2_NMU128_DATA_SZ 32

// Attribute addresses
//

`define NOC2_NMU128__REG_ADDR_DST0    32'h00000000
`define NOC2_NMU128__REG_ADDR_DST0_SZ 18

`define NOC2_NMU128__REG_ADDR_DST1    32'h00000001
`define NOC2_NMU128__REG_ADDR_DST1_SZ 18

`define NOC2_NMU128__REG_ADDR_DST10    32'h00000002
`define NOC2_NMU128__REG_ADDR_DST10_SZ 18

`define NOC2_NMU128__REG_ADDR_DST11    32'h00000003
`define NOC2_NMU128__REG_ADDR_DST11_SZ 18

`define NOC2_NMU128__REG_ADDR_DST12    32'h00000004
`define NOC2_NMU128__REG_ADDR_DST12_SZ 18

`define NOC2_NMU128__REG_ADDR_DST13    32'h00000005
`define NOC2_NMU128__REG_ADDR_DST13_SZ 18

`define NOC2_NMU128__REG_ADDR_DST14    32'h00000006
`define NOC2_NMU128__REG_ADDR_DST14_SZ 18

`define NOC2_NMU128__REG_ADDR_DST15    32'h00000007
`define NOC2_NMU128__REG_ADDR_DST15_SZ 18

`define NOC2_NMU128__REG_ADDR_DST16    32'h00000008
`define NOC2_NMU128__REG_ADDR_DST16_SZ 18

`define NOC2_NMU128__REG_ADDR_DST17    32'h00000009
`define NOC2_NMU128__REG_ADDR_DST17_SZ 18

`define NOC2_NMU128__REG_ADDR_DST18    32'h0000000a
`define NOC2_NMU128__REG_ADDR_DST18_SZ 18

`define NOC2_NMU128__REG_ADDR_DST19    32'h0000000b
`define NOC2_NMU128__REG_ADDR_DST19_SZ 18

`define NOC2_NMU128__REG_ADDR_DST2    32'h0000000c
`define NOC2_NMU128__REG_ADDR_DST2_SZ 18

`define NOC2_NMU128__REG_ADDR_DST20    32'h0000000d
`define NOC2_NMU128__REG_ADDR_DST20_SZ 18

`define NOC2_NMU128__REG_ADDR_DST21    32'h0000000e
`define NOC2_NMU128__REG_ADDR_DST21_SZ 18

`define NOC2_NMU128__REG_ADDR_DST22    32'h0000000f
`define NOC2_NMU128__REG_ADDR_DST22_SZ 18

`define NOC2_NMU128__REG_ADDR_DST23    32'h00000010
`define NOC2_NMU128__REG_ADDR_DST23_SZ 18

`define NOC2_NMU128__REG_ADDR_DST24    32'h00000011
`define NOC2_NMU128__REG_ADDR_DST24_SZ 18

`define NOC2_NMU128__REG_ADDR_DST25    32'h00000012
`define NOC2_NMU128__REG_ADDR_DST25_SZ 18

`define NOC2_NMU128__REG_ADDR_DST26    32'h00000013
`define NOC2_NMU128__REG_ADDR_DST26_SZ 18

`define NOC2_NMU128__REG_ADDR_DST27    32'h00000014
`define NOC2_NMU128__REG_ADDR_DST27_SZ 18

`define NOC2_NMU128__REG_ADDR_DST28    32'h00000015
`define NOC2_NMU128__REG_ADDR_DST28_SZ 18

`define NOC2_NMU128__REG_ADDR_DST29    32'h00000016
`define NOC2_NMU128__REG_ADDR_DST29_SZ 18

`define NOC2_NMU128__REG_ADDR_DST3    32'h00000017
`define NOC2_NMU128__REG_ADDR_DST3_SZ 18

`define NOC2_NMU128__REG_ADDR_DST30    32'h00000018
`define NOC2_NMU128__REG_ADDR_DST30_SZ 18

`define NOC2_NMU128__REG_ADDR_DST31    32'h00000019
`define NOC2_NMU128__REG_ADDR_DST31_SZ 18

`define NOC2_NMU128__REG_ADDR_DST4    32'h0000001a
`define NOC2_NMU128__REG_ADDR_DST4_SZ 18

`define NOC2_NMU128__REG_ADDR_DST5    32'h0000001b
`define NOC2_NMU128__REG_ADDR_DST5_SZ 18

`define NOC2_NMU128__REG_ADDR_DST6    32'h0000001c
`define NOC2_NMU128__REG_ADDR_DST6_SZ 18

`define NOC2_NMU128__REG_ADDR_DST7    32'h0000001d
`define NOC2_NMU128__REG_ADDR_DST7_SZ 18

`define NOC2_NMU128__REG_ADDR_DST8    32'h0000001e
`define NOC2_NMU128__REG_ADDR_DST8_SZ 18

`define NOC2_NMU128__REG_ADDR_DST9    32'h0000001f
`define NOC2_NMU128__REG_ADDR_DST9_SZ 18

`define NOC2_NMU128__REG_ADDR_ENABLE    32'h00000020
`define NOC2_NMU128__REG_ADDR_ENABLE_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR0    32'h00000021
`define NOC2_NMU128__REG_ADDR_MADDR0_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR1    32'h00000022
`define NOC2_NMU128__REG_ADDR_MADDR1_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR10    32'h00000023
`define NOC2_NMU128__REG_ADDR_MADDR10_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR11    32'h00000024
`define NOC2_NMU128__REG_ADDR_MADDR11_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR12    32'h00000025
`define NOC2_NMU128__REG_ADDR_MADDR12_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR13    32'h00000026
`define NOC2_NMU128__REG_ADDR_MADDR13_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR14    32'h00000027
`define NOC2_NMU128__REG_ADDR_MADDR14_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR15    32'h00000028
`define NOC2_NMU128__REG_ADDR_MADDR15_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR16    32'h00000029
`define NOC2_NMU128__REG_ADDR_MADDR16_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR17    32'h0000002a
`define NOC2_NMU128__REG_ADDR_MADDR17_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR18    32'h0000002b
`define NOC2_NMU128__REG_ADDR_MADDR18_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR19    32'h0000002c
`define NOC2_NMU128__REG_ADDR_MADDR19_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR2    32'h0000002d
`define NOC2_NMU128__REG_ADDR_MADDR2_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR20    32'h0000002e
`define NOC2_NMU128__REG_ADDR_MADDR20_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR21    32'h0000002f
`define NOC2_NMU128__REG_ADDR_MADDR21_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR22    32'h00000030
`define NOC2_NMU128__REG_ADDR_MADDR22_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR23    32'h00000031
`define NOC2_NMU128__REG_ADDR_MADDR23_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR24    32'h00000032
`define NOC2_NMU128__REG_ADDR_MADDR24_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR25    32'h00000033
`define NOC2_NMU128__REG_ADDR_MADDR25_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR26    32'h00000034
`define NOC2_NMU128__REG_ADDR_MADDR26_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR27    32'h00000035
`define NOC2_NMU128__REG_ADDR_MADDR27_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR28    32'h00000036
`define NOC2_NMU128__REG_ADDR_MADDR28_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR29    32'h00000037
`define NOC2_NMU128__REG_ADDR_MADDR29_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR3    32'h00000038
`define NOC2_NMU128__REG_ADDR_MADDR3_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR30    32'h00000039
`define NOC2_NMU128__REG_ADDR_MADDR30_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR31    32'h0000003a
`define NOC2_NMU128__REG_ADDR_MADDR31_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR4    32'h0000003b
`define NOC2_NMU128__REG_ADDR_MADDR4_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR5    32'h0000003c
`define NOC2_NMU128__REG_ADDR_MADDR5_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR6    32'h0000003d
`define NOC2_NMU128__REG_ADDR_MADDR6_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR7    32'h0000003e
`define NOC2_NMU128__REG_ADDR_MADDR7_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR8    32'h0000003f
`define NOC2_NMU128__REG_ADDR_MADDR8_SZ 32

`define NOC2_NMU128__REG_ADDR_MADDR9    32'h00000040
`define NOC2_NMU128__REG_ADDR_MADDR9_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK0    32'h00000041
`define NOC2_NMU128__REG_ADDR_MASK0_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK1    32'h00000042
`define NOC2_NMU128__REG_ADDR_MASK1_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK10    32'h00000043
`define NOC2_NMU128__REG_ADDR_MASK10_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK11    32'h00000044
`define NOC2_NMU128__REG_ADDR_MASK11_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK12    32'h00000045
`define NOC2_NMU128__REG_ADDR_MASK12_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK13    32'h00000046
`define NOC2_NMU128__REG_ADDR_MASK13_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK14    32'h00000047
`define NOC2_NMU128__REG_ADDR_MASK14_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK15    32'h00000048
`define NOC2_NMU128__REG_ADDR_MASK15_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK16    32'h00000049
`define NOC2_NMU128__REG_ADDR_MASK16_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK17    32'h0000004a
`define NOC2_NMU128__REG_ADDR_MASK17_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK18    32'h0000004b
`define NOC2_NMU128__REG_ADDR_MASK18_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK19    32'h0000004c
`define NOC2_NMU128__REG_ADDR_MASK19_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK2    32'h0000004d
`define NOC2_NMU128__REG_ADDR_MASK2_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK20    32'h0000004e
`define NOC2_NMU128__REG_ADDR_MASK20_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK21    32'h0000004f
`define NOC2_NMU128__REG_ADDR_MASK21_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK22    32'h00000050
`define NOC2_NMU128__REG_ADDR_MASK22_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK23    32'h00000051
`define NOC2_NMU128__REG_ADDR_MASK23_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK24    32'h00000052
`define NOC2_NMU128__REG_ADDR_MASK24_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK25    32'h00000053
`define NOC2_NMU128__REG_ADDR_MASK25_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK26    32'h00000054
`define NOC2_NMU128__REG_ADDR_MASK26_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK27    32'h00000055
`define NOC2_NMU128__REG_ADDR_MASK27_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK28    32'h00000056
`define NOC2_NMU128__REG_ADDR_MASK28_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK29    32'h00000057
`define NOC2_NMU128__REG_ADDR_MASK29_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK3    32'h00000058
`define NOC2_NMU128__REG_ADDR_MASK3_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK30    32'h00000059
`define NOC2_NMU128__REG_ADDR_MASK30_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK31    32'h0000005a
`define NOC2_NMU128__REG_ADDR_MASK31_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK4    32'h0000005b
`define NOC2_NMU128__REG_ADDR_MASK4_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK5    32'h0000005c
`define NOC2_NMU128__REG_ADDR_MASK5_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK6    32'h0000005d
`define NOC2_NMU128__REG_ADDR_MASK6_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK7    32'h0000005e
`define NOC2_NMU128__REG_ADDR_MASK7_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK8    32'h0000005f
`define NOC2_NMU128__REG_ADDR_MASK8_SZ 32

`define NOC2_NMU128__REG_ADDR_MASK9    32'h00000060
`define NOC2_NMU128__REG_ADDR_MASK9_SZ 32

`define NOC2_NMU128__REG_ADDR_REMAP    32'h00000061
`define NOC2_NMU128__REG_ADDR_REMAP_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR0    32'h00000062
`define NOC2_NMU128__REG_ADDR_RPADDR0_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR1    32'h00000063
`define NOC2_NMU128__REG_ADDR_RPADDR1_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR10    32'h00000064
`define NOC2_NMU128__REG_ADDR_RPADDR10_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR11    32'h00000065
`define NOC2_NMU128__REG_ADDR_RPADDR11_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR12    32'h00000066
`define NOC2_NMU128__REG_ADDR_RPADDR12_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR13    32'h00000067
`define NOC2_NMU128__REG_ADDR_RPADDR13_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR14    32'h00000068
`define NOC2_NMU128__REG_ADDR_RPADDR14_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR15    32'h00000069
`define NOC2_NMU128__REG_ADDR_RPADDR15_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR16    32'h0000006a
`define NOC2_NMU128__REG_ADDR_RPADDR16_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR17    32'h0000006b
`define NOC2_NMU128__REG_ADDR_RPADDR17_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR18    32'h0000006c
`define NOC2_NMU128__REG_ADDR_RPADDR18_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR19    32'h0000006d
`define NOC2_NMU128__REG_ADDR_RPADDR19_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR2    32'h0000006e
`define NOC2_NMU128__REG_ADDR_RPADDR2_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR20    32'h0000006f
`define NOC2_NMU128__REG_ADDR_RPADDR20_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR21    32'h00000070
`define NOC2_NMU128__REG_ADDR_RPADDR21_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR22    32'h00000071
`define NOC2_NMU128__REG_ADDR_RPADDR22_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR23    32'h00000072
`define NOC2_NMU128__REG_ADDR_RPADDR23_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR24    32'h00000073
`define NOC2_NMU128__REG_ADDR_RPADDR24_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR25    32'h00000074
`define NOC2_NMU128__REG_ADDR_RPADDR25_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR26    32'h00000075
`define NOC2_NMU128__REG_ADDR_RPADDR26_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR27    32'h00000076
`define NOC2_NMU128__REG_ADDR_RPADDR27_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR28    32'h00000077
`define NOC2_NMU128__REG_ADDR_RPADDR28_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR29    32'h00000078
`define NOC2_NMU128__REG_ADDR_RPADDR29_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR3    32'h00000079
`define NOC2_NMU128__REG_ADDR_RPADDR3_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR30    32'h0000007a
`define NOC2_NMU128__REG_ADDR_RPADDR30_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR31    32'h0000007b
`define NOC2_NMU128__REG_ADDR_RPADDR31_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR4    32'h0000007c
`define NOC2_NMU128__REG_ADDR_RPADDR4_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR5    32'h0000007d
`define NOC2_NMU128__REG_ADDR_RPADDR5_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR6    32'h0000007e
`define NOC2_NMU128__REG_ADDR_RPADDR6_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR7    32'h0000007f
`define NOC2_NMU128__REG_ADDR_RPADDR7_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR8    32'h00000080
`define NOC2_NMU128__REG_ADDR_RPADDR8_SZ 32

`define NOC2_NMU128__REG_ADDR_RPADDR9    32'h00000081
`define NOC2_NMU128__REG_ADDR_RPADDR9_SZ 32

`define NOC2_NMU128__REG_ADR_MAP_CPM    32'h00000082
`define NOC2_NMU128__REG_ADR_MAP_CPM_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_FPD_AFI_FS_0    32'h00000083
`define NOC2_NMU128__REG_ADR_MAP_FPD_AFI_FS_0_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_FPD_AFI_FS_1    32'h00000084
`define NOC2_NMU128__REG_ADR_MAP_FPD_AFI_FS_1_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_FPD_GIC    32'h00000085
`define NOC2_NMU128__REG_ADR_MAP_FPD_GIC_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_HNIC    32'h00000086
`define NOC2_NMU128__REG_ADR_MAP_HNIC_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_LPD_AFI_FS    32'h00000087
`define NOC2_NMU128__REG_ADR_MAP_LPD_AFI_FS_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_0    32'h00000088
`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_0_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_1    32'h00000089
`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_1_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_2    32'h0000008a
`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_2_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_3    32'h0000008b
`define NOC2_NMU128__REG_ADR_MAP_ME_ARRAY_3_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_OCM    32'h0000008c
`define NOC2_NMU128__REG_ADR_MAP_OCM_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PCIE    32'h0000008d
`define NOC2_NMU128__REG_ADR_MAP_PCIE_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PMC    32'h0000008e
`define NOC2_NMU128__REG_ADR_MAP_PMC_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_0    32'h0000008f
`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_0_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_1    32'h00000090
`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_1_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_2    32'h00000091
`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_2_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_3    32'h00000092
`define NOC2_NMU128__REG_ADR_MAP_PMC_ALIAS_3_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_XPDS    32'h00000093
`define NOC2_NMU128__REG_ADR_MAP_XPDS_SZ 15

`define NOC2_NMU128__REG_ADR_MAP_XSPI    32'h00000094
`define NOC2_NMU128__REG_ADR_MAP_XSPI_SZ 15

`define NOC2_NMU128__REG_AFWS_EN    32'h00000095
`define NOC2_NMU128__REG_AFWS_EN_SZ 1

`define NOC2_NMU128__REG_AFWS_INTR_EN    32'h00000096
`define NOC2_NMU128__REG_AFWS_INTR_EN_SZ 1

`define NOC2_NMU128__REG_AFWS_TIMEOUT_ERR_EN    32'h00000097
`define NOC2_NMU128__REG_AFWS_TIMEOUT_ERR_EN_SZ 4

`define NOC2_NMU128__REG_AXI_NON_MOD_DISABLE    32'h00000098
`define NOC2_NMU128__REG_AXI_NON_MOD_DISABLE_SZ 1

`define NOC2_NMU128__REG_AXI_PAR_CHK    32'h00000099
`define NOC2_NMU128__REG_AXI_PAR_CHK_SZ 2

`define NOC2_NMU128__REG_CHOPSIZE    32'h0000009a
`define NOC2_NMU128__REG_CHOPSIZE_SZ 4

`define NOC2_NMU128__REG_DDR_ADR_MAP0_0    32'h0000009b
`define NOC2_NMU128__REG_DDR_ADR_MAP0_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP0_1    32'h0000009c
`define NOC2_NMU128__REG_DDR_ADR_MAP0_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP1_0    32'h0000009d
`define NOC2_NMU128__REG_DDR_ADR_MAP1_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP1_1    32'h0000009e
`define NOC2_NMU128__REG_DDR_ADR_MAP1_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP2_0    32'h0000009f
`define NOC2_NMU128__REG_DDR_ADR_MAP2_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP2_1    32'h000000a0
`define NOC2_NMU128__REG_DDR_ADR_MAP2_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP3_0    32'h000000a1
`define NOC2_NMU128__REG_DDR_ADR_MAP3_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP3_1    32'h000000a2
`define NOC2_NMU128__REG_DDR_ADR_MAP3_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP4_0    32'h000000a3
`define NOC2_NMU128__REG_DDR_ADR_MAP4_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP4_1    32'h000000a4
`define NOC2_NMU128__REG_DDR_ADR_MAP4_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP5_0    32'h000000a5
`define NOC2_NMU128__REG_DDR_ADR_MAP5_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP5_1    32'h000000a6
`define NOC2_NMU128__REG_DDR_ADR_MAP5_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP6_0    32'h000000a7
`define NOC2_NMU128__REG_DDR_ADR_MAP6_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP6_1    32'h000000a8
`define NOC2_NMU128__REG_DDR_ADR_MAP6_1_SZ 6

`define NOC2_NMU128__REG_DDR_ADR_MAP7_0    32'h000000a9
`define NOC2_NMU128__REG_DDR_ADR_MAP7_0_SZ 32

`define NOC2_NMU128__REG_DDR_ADR_MAP7_1    32'h000000aa
`define NOC2_NMU128__REG_DDR_ADR_MAP7_1_SZ 6

`define NOC2_NMU128__REG_DDR_DST_MAP0    32'h000000ab
`define NOC2_NMU128__REG_DDR_DST_MAP0_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP1    32'h000000ac
`define NOC2_NMU128__REG_DDR_DST_MAP1_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP10    32'h000000ad
`define NOC2_NMU128__REG_DDR_DST_MAP10_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP11    32'h000000ae
`define NOC2_NMU128__REG_DDR_DST_MAP11_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP12    32'h000000af
`define NOC2_NMU128__REG_DDR_DST_MAP12_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP13    32'h000000b0
`define NOC2_NMU128__REG_DDR_DST_MAP13_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP14    32'h000000b1
`define NOC2_NMU128__REG_DDR_DST_MAP14_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP15    32'h000000b2
`define NOC2_NMU128__REG_DDR_DST_MAP15_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP2    32'h000000b3
`define NOC2_NMU128__REG_DDR_DST_MAP2_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP3    32'h000000b4
`define NOC2_NMU128__REG_DDR_DST_MAP3_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP4    32'h000000b5
`define NOC2_NMU128__REG_DDR_DST_MAP4_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP5    32'h000000b6
`define NOC2_NMU128__REG_DDR_DST_MAP5_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP6    32'h000000b7
`define NOC2_NMU128__REG_DDR_DST_MAP6_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP7    32'h000000b8
`define NOC2_NMU128__REG_DDR_DST_MAP7_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP8    32'h000000b9
`define NOC2_NMU128__REG_DDR_DST_MAP8_SZ 12

`define NOC2_NMU128__REG_DDR_DST_MAP9    32'h000000ba
`define NOC2_NMU128__REG_DDR_DST_MAP9_SZ 12

`define NOC2_NMU128__REG_DWIDTH    32'h000000bb
`define NOC2_NMU128__REG_DWIDTH_SZ 3

`define NOC2_NMU128__REG_ECC_CHK_EN    32'h000000bc
`define NOC2_NMU128__REG_ECC_CHK_EN_SZ 1

`define NOC2_NMU128__REG_HBM_MAP_T0_CH0    32'h000000bd
`define NOC2_NMU128__REG_HBM_MAP_T0_CH0_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH1    32'h000000be
`define NOC2_NMU128__REG_HBM_MAP_T0_CH1_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH10    32'h000000bf
`define NOC2_NMU128__REG_HBM_MAP_T0_CH10_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH11    32'h000000c0
`define NOC2_NMU128__REG_HBM_MAP_T0_CH11_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH12    32'h000000c1
`define NOC2_NMU128__REG_HBM_MAP_T0_CH12_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH13    32'h000000c2
`define NOC2_NMU128__REG_HBM_MAP_T0_CH13_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH14    32'h000000c3
`define NOC2_NMU128__REG_HBM_MAP_T0_CH14_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH15    32'h000000c4
`define NOC2_NMU128__REG_HBM_MAP_T0_CH15_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH2    32'h000000c5
`define NOC2_NMU128__REG_HBM_MAP_T0_CH2_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH3    32'h000000c6
`define NOC2_NMU128__REG_HBM_MAP_T0_CH3_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH4    32'h000000c7
`define NOC2_NMU128__REG_HBM_MAP_T0_CH4_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH5    32'h000000c8
`define NOC2_NMU128__REG_HBM_MAP_T0_CH5_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH6    32'h000000c9
`define NOC2_NMU128__REG_HBM_MAP_T0_CH6_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH7    32'h000000ca
`define NOC2_NMU128__REG_HBM_MAP_T0_CH7_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH8    32'h000000cb
`define NOC2_NMU128__REG_HBM_MAP_T0_CH8_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T0_CH9    32'h000000cc
`define NOC2_NMU128__REG_HBM_MAP_T0_CH9_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH0    32'h000000cd
`define NOC2_NMU128__REG_HBM_MAP_T1_CH0_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH1    32'h000000ce
`define NOC2_NMU128__REG_HBM_MAP_T1_CH1_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH10    32'h000000cf
`define NOC2_NMU128__REG_HBM_MAP_T1_CH10_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH11    32'h000000d0
`define NOC2_NMU128__REG_HBM_MAP_T1_CH11_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH12    32'h000000d1
`define NOC2_NMU128__REG_HBM_MAP_T1_CH12_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH13    32'h000000d2
`define NOC2_NMU128__REG_HBM_MAP_T1_CH13_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH14    32'h000000d3
`define NOC2_NMU128__REG_HBM_MAP_T1_CH14_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH15    32'h000000d4
`define NOC2_NMU128__REG_HBM_MAP_T1_CH15_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH2    32'h000000d5
`define NOC2_NMU128__REG_HBM_MAP_T1_CH2_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH3    32'h000000d6
`define NOC2_NMU128__REG_HBM_MAP_T1_CH3_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH4    32'h000000d7
`define NOC2_NMU128__REG_HBM_MAP_T1_CH4_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH5    32'h000000d8
`define NOC2_NMU128__REG_HBM_MAP_T1_CH5_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH6    32'h000000d9
`define NOC2_NMU128__REG_HBM_MAP_T1_CH6_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH7    32'h000000da
`define NOC2_NMU128__REG_HBM_MAP_T1_CH7_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH8    32'h000000db
`define NOC2_NMU128__REG_HBM_MAP_T1_CH8_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T1_CH9    32'h000000dc
`define NOC2_NMU128__REG_HBM_MAP_T1_CH9_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH0    32'h000000dd
`define NOC2_NMU128__REG_HBM_MAP_T2_CH0_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH1    32'h000000de
`define NOC2_NMU128__REG_HBM_MAP_T2_CH1_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH10    32'h000000df
`define NOC2_NMU128__REG_HBM_MAP_T2_CH10_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH11    32'h000000e0
`define NOC2_NMU128__REG_HBM_MAP_T2_CH11_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH12    32'h000000e1
`define NOC2_NMU128__REG_HBM_MAP_T2_CH12_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH13    32'h000000e2
`define NOC2_NMU128__REG_HBM_MAP_T2_CH13_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH14    32'h000000e3
`define NOC2_NMU128__REG_HBM_MAP_T2_CH14_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH15    32'h000000e4
`define NOC2_NMU128__REG_HBM_MAP_T2_CH15_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH2    32'h000000e5
`define NOC2_NMU128__REG_HBM_MAP_T2_CH2_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH3    32'h000000e6
`define NOC2_NMU128__REG_HBM_MAP_T2_CH3_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH4    32'h000000e7
`define NOC2_NMU128__REG_HBM_MAP_T2_CH4_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH5    32'h000000e8
`define NOC2_NMU128__REG_HBM_MAP_T2_CH5_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH6    32'h000000e9
`define NOC2_NMU128__REG_HBM_MAP_T2_CH6_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH7    32'h000000ea
`define NOC2_NMU128__REG_HBM_MAP_T2_CH7_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH8    32'h000000eb
`define NOC2_NMU128__REG_HBM_MAP_T2_CH8_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T2_CH9    32'h000000ec
`define NOC2_NMU128__REG_HBM_MAP_T2_CH9_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH0    32'h000000ed
`define NOC2_NMU128__REG_HBM_MAP_T3_CH0_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH1    32'h000000ee
`define NOC2_NMU128__REG_HBM_MAP_T3_CH1_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH10    32'h000000ef
`define NOC2_NMU128__REG_HBM_MAP_T3_CH10_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH11    32'h000000f0
`define NOC2_NMU128__REG_HBM_MAP_T3_CH11_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH12    32'h000000f1
`define NOC2_NMU128__REG_HBM_MAP_T3_CH12_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH13    32'h000000f2
`define NOC2_NMU128__REG_HBM_MAP_T3_CH13_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH14    32'h000000f3
`define NOC2_NMU128__REG_HBM_MAP_T3_CH14_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH15    32'h000000f4
`define NOC2_NMU128__REG_HBM_MAP_T3_CH15_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH2    32'h000000f5
`define NOC2_NMU128__REG_HBM_MAP_T3_CH2_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH3    32'h000000f6
`define NOC2_NMU128__REG_HBM_MAP_T3_CH3_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH4    32'h000000f7
`define NOC2_NMU128__REG_HBM_MAP_T3_CH4_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH5    32'h000000f8
`define NOC2_NMU128__REG_HBM_MAP_T3_CH5_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH6    32'h000000f9
`define NOC2_NMU128__REG_HBM_MAP_T3_CH6_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH7    32'h000000fa
`define NOC2_NMU128__REG_HBM_MAP_T3_CH7_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH8    32'h000000fb
`define NOC2_NMU128__REG_HBM_MAP_T3_CH8_SZ 15

`define NOC2_NMU128__REG_HBM_MAP_T3_CH9    32'h000000fc
`define NOC2_NMU128__REG_HBM_MAP_T3_CH9_SZ 15

`define NOC2_NMU128__REG_MODE_SELECT    32'h000000fd
`define NOC2_NMU128__REG_MODE_SELECT_SZ 16

`define NOC2_NMU128__REG_NMU_BYPASS_EN    32'h000000fe
`define NOC2_NMU128__REG_NMU_BYPASS_EN_SZ 1

`define NOC2_NMU128__REG_OUTSTANDING_RD_TXN    32'h000000ff
`define NOC2_NMU128__REG_OUTSTANDING_RD_TXN_SZ 7

`define NOC2_NMU128__REG_OUTSTANDING_WR_TXN    32'h00000100
`define NOC2_NMU128__REG_OUTSTANDING_WR_TXN_SZ 7

`define NOC2_NMU128__REG_PRIORITY    32'h00000101
`define NOC2_NMU128__REG_PRIORITY_SZ 2

`define NOC2_NMU128__REG_RD_AXPROT_SEL    32'h00000102
`define NOC2_NMU128__REG_RD_AXPROT_SEL_SZ 6

`define NOC2_NMU128__REG_RD_RATE_CREDIT_DROP    32'h00000103
`define NOC2_NMU128__REG_RD_RATE_CREDIT_DROP_SZ 10

`define NOC2_NMU128__REG_RD_RATE_CREDIT_LIMIT    32'h00000104
`define NOC2_NMU128__REG_RD_RATE_CREDIT_LIMIT_SZ 14

`define NOC2_NMU128__REG_RD_VCA_TOKEN0    32'h00000105
`define NOC2_NMU128__REG_RD_VCA_TOKEN0_SZ 8

`define NOC2_NMU128__REG_RESP_SRC_ID_MASK    32'h00000106
`define NOC2_NMU128__REG_RESP_SRC_ID_MASK_SZ 12

`define NOC2_NMU128__REG_RPOISON_TO_SLVERR    32'h00000107
`define NOC2_NMU128__REG_RPOISON_TO_SLVERR_SZ 1

`define NOC2_NMU128__REG_RROB_RAM_SETTING    32'h00000108
`define NOC2_NMU128__REG_RROB_RAM_SETTING_SZ 9

`define NOC2_NMU128__REG_SMID_SEL    32'h00000109
`define NOC2_NMU128__REG_SMID_SEL_SZ 20

`define NOC2_NMU128__REG_SRC    32'h0000010a
`define NOC2_NMU128__REG_SRC_SZ 12

`define NOC2_NMU128__REG_TBASE_AXI_TIMEOUT    32'h0000010b
`define NOC2_NMU128__REG_TBASE_AXI_TIMEOUT_SZ 4

`define NOC2_NMU128__REG_TBASE_MODE_RLIMIT_RD    32'h0000010c
`define NOC2_NMU128__REG_TBASE_MODE_RLIMIT_RD_SZ 3

`define NOC2_NMU128__REG_TBASE_MODE_RLIMIT_WR    32'h0000010d
`define NOC2_NMU128__REG_TBASE_MODE_RLIMIT_WR_SZ 3

`define NOC2_NMU128__REG_TBASE_TRK_TIMEOUT    32'h0000010e
`define NOC2_NMU128__REG_TBASE_TRK_TIMEOUT_SZ 4

`define NOC2_NMU128__REG_USER_DST0    32'h0000010f
`define NOC2_NMU128__REG_USER_DST0_SZ 15

`define NOC2_NMU128__REG_USER_DST1    32'h00000110
`define NOC2_NMU128__REG_USER_DST1_SZ 15

`define NOC2_NMU128__REG_USER_DST10    32'h00000111
`define NOC2_NMU128__REG_USER_DST10_SZ 15

`define NOC2_NMU128__REG_USER_DST11    32'h00000112
`define NOC2_NMU128__REG_USER_DST11_SZ 15

`define NOC2_NMU128__REG_USER_DST12    32'h00000113
`define NOC2_NMU128__REG_USER_DST12_SZ 15

`define NOC2_NMU128__REG_USER_DST13    32'h00000114
`define NOC2_NMU128__REG_USER_DST13_SZ 15

`define NOC2_NMU128__REG_USER_DST14    32'h00000115
`define NOC2_NMU128__REG_USER_DST14_SZ 15

`define NOC2_NMU128__REG_USER_DST15    32'h00000116
`define NOC2_NMU128__REG_USER_DST15_SZ 15

`define NOC2_NMU128__REG_USER_DST2    32'h00000117
`define NOC2_NMU128__REG_USER_DST2_SZ 15

`define NOC2_NMU128__REG_USER_DST3    32'h00000118
`define NOC2_NMU128__REG_USER_DST3_SZ 15

`define NOC2_NMU128__REG_USER_DST4    32'h00000119
`define NOC2_NMU128__REG_USER_DST4_SZ 15

`define NOC2_NMU128__REG_USER_DST5    32'h0000011a
`define NOC2_NMU128__REG_USER_DST5_SZ 15

`define NOC2_NMU128__REG_USER_DST6    32'h0000011b
`define NOC2_NMU128__REG_USER_DST6_SZ 15

`define NOC2_NMU128__REG_USER_DST7    32'h0000011c
`define NOC2_NMU128__REG_USER_DST7_SZ 15

`define NOC2_NMU128__REG_USER_DST8    32'h0000011d
`define NOC2_NMU128__REG_USER_DST8_SZ 15

`define NOC2_NMU128__REG_USER_DST9    32'h0000011e
`define NOC2_NMU128__REG_USER_DST9_SZ 15

`define NOC2_NMU128__REG_USER_REMAP_CTRL    32'h0000011f
`define NOC2_NMU128__REG_USER_REMAP_CTRL_SZ 1

`define NOC2_NMU128__REG_VC_MAP    32'h00000120
`define NOC2_NMU128__REG_VC_MAP_SZ 12

`define NOC2_NMU128__REG_WBUF_LAUNCH_SIZE    32'h00000121
`define NOC2_NMU128__REG_WBUF_LAUNCH_SIZE_SZ 6

`define NOC2_NMU128__REG_WBUF_RAM_SETTING    32'h00000122
`define NOC2_NMU128__REG_WBUF_RAM_SETTING_SZ 9

`define NOC2_NMU128__REG_WR_AXPROT_SEL    32'h00000123
`define NOC2_NMU128__REG_WR_AXPROT_SEL_SZ 6

`define NOC2_NMU128__REG_WR_RATE_CREDIT_DROP    32'h00000124
`define NOC2_NMU128__REG_WR_RATE_CREDIT_DROP_SZ 10

`define NOC2_NMU128__REG_WR_RATE_CREDIT_LIMIT    32'h00000125
`define NOC2_NMU128__REG_WR_RATE_CREDIT_LIMIT_SZ 14

`define NOC2_NMU128__REG_WR_VCA_TOKEN0    32'h00000126
`define NOC2_NMU128__REG_WR_VCA_TOKEN0_SZ 8

`endif  // B_NOC2_NMU128_DEFINES_VH