// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC_NMU128_DEFINES_VH
`else
`define B_NOC_NMU128_DEFINES_VH

// Look-up table parameters
//

`define NOC_NMU128_ADDR_N  190
`define NOC_NMU128_ADDR_SZ 32
`define NOC_NMU128_DATA_SZ 32

// Attribute addresses
//

`define NOC_NMU128__REG_ADDR_DST0    32'h00000000
`define NOC_NMU128__REG_ADDR_DST0_SZ 16

`define NOC_NMU128__REG_ADDR_DST1    32'h00000001
`define NOC_NMU128__REG_ADDR_DST1_SZ 16

`define NOC_NMU128__REG_ADDR_DST10    32'h00000002
`define NOC_NMU128__REG_ADDR_DST10_SZ 16

`define NOC_NMU128__REG_ADDR_DST11    32'h00000003
`define NOC_NMU128__REG_ADDR_DST11_SZ 16

`define NOC_NMU128__REG_ADDR_DST12    32'h00000004
`define NOC_NMU128__REG_ADDR_DST12_SZ 16

`define NOC_NMU128__REG_ADDR_DST13    32'h00000005
`define NOC_NMU128__REG_ADDR_DST13_SZ 16

`define NOC_NMU128__REG_ADDR_DST14    32'h00000006
`define NOC_NMU128__REG_ADDR_DST14_SZ 16

`define NOC_NMU128__REG_ADDR_DST15    32'h00000007
`define NOC_NMU128__REG_ADDR_DST15_SZ 16

`define NOC_NMU128__REG_ADDR_DST2    32'h00000008
`define NOC_NMU128__REG_ADDR_DST2_SZ 16

`define NOC_NMU128__REG_ADDR_DST3    32'h00000009
`define NOC_NMU128__REG_ADDR_DST3_SZ 16

`define NOC_NMU128__REG_ADDR_DST4    32'h0000000a
`define NOC_NMU128__REG_ADDR_DST4_SZ 16

`define NOC_NMU128__REG_ADDR_DST5    32'h0000000b
`define NOC_NMU128__REG_ADDR_DST5_SZ 16

`define NOC_NMU128__REG_ADDR_DST6    32'h0000000c
`define NOC_NMU128__REG_ADDR_DST6_SZ 16

`define NOC_NMU128__REG_ADDR_DST7    32'h0000000d
`define NOC_NMU128__REG_ADDR_DST7_SZ 16

`define NOC_NMU128__REG_ADDR_DST8    32'h0000000e
`define NOC_NMU128__REG_ADDR_DST8_SZ 16

`define NOC_NMU128__REG_ADDR_DST9    32'h0000000f
`define NOC_NMU128__REG_ADDR_DST9_SZ 16

`define NOC_NMU128__REG_ADDR_ENABLE    32'h00000010
`define NOC_NMU128__REG_ADDR_ENABLE_SZ 16

`define NOC_NMU128__REG_ADDR_MADDR0    32'h00000011
`define NOC_NMU128__REG_ADDR_MADDR0_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR1    32'h00000012
`define NOC_NMU128__REG_ADDR_MADDR1_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR10    32'h00000013
`define NOC_NMU128__REG_ADDR_MADDR10_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR11    32'h00000014
`define NOC_NMU128__REG_ADDR_MADDR11_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR12    32'h00000015
`define NOC_NMU128__REG_ADDR_MADDR12_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR13    32'h00000016
`define NOC_NMU128__REG_ADDR_MADDR13_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR14    32'h00000017
`define NOC_NMU128__REG_ADDR_MADDR14_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR15    32'h00000018
`define NOC_NMU128__REG_ADDR_MADDR15_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR2    32'h00000019
`define NOC_NMU128__REG_ADDR_MADDR2_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR3    32'h0000001a
`define NOC_NMU128__REG_ADDR_MADDR3_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR4    32'h0000001b
`define NOC_NMU128__REG_ADDR_MADDR4_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR5    32'h0000001c
`define NOC_NMU128__REG_ADDR_MADDR5_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR6    32'h0000001d
`define NOC_NMU128__REG_ADDR_MADDR6_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR7    32'h0000001e
`define NOC_NMU128__REG_ADDR_MADDR7_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR8    32'h0000001f
`define NOC_NMU128__REG_ADDR_MADDR8_SZ 32

`define NOC_NMU128__REG_ADDR_MADDR9    32'h00000020
`define NOC_NMU128__REG_ADDR_MADDR9_SZ 32

`define NOC_NMU128__REG_ADDR_MASK0    32'h00000021
`define NOC_NMU128__REG_ADDR_MASK0_SZ 32

`define NOC_NMU128__REG_ADDR_MASK1    32'h00000022
`define NOC_NMU128__REG_ADDR_MASK1_SZ 32

`define NOC_NMU128__REG_ADDR_MASK10    32'h00000023
`define NOC_NMU128__REG_ADDR_MASK10_SZ 32

`define NOC_NMU128__REG_ADDR_MASK11    32'h00000024
`define NOC_NMU128__REG_ADDR_MASK11_SZ 32

`define NOC_NMU128__REG_ADDR_MASK12    32'h00000025
`define NOC_NMU128__REG_ADDR_MASK12_SZ 32

`define NOC_NMU128__REG_ADDR_MASK13    32'h00000026
`define NOC_NMU128__REG_ADDR_MASK13_SZ 32

`define NOC_NMU128__REG_ADDR_MASK14    32'h00000027
`define NOC_NMU128__REG_ADDR_MASK14_SZ 32

`define NOC_NMU128__REG_ADDR_MASK15    32'h00000028
`define NOC_NMU128__REG_ADDR_MASK15_SZ 32

`define NOC_NMU128__REG_ADDR_MASK2    32'h00000029
`define NOC_NMU128__REG_ADDR_MASK2_SZ 32

`define NOC_NMU128__REG_ADDR_MASK3    32'h0000002a
`define NOC_NMU128__REG_ADDR_MASK3_SZ 32

`define NOC_NMU128__REG_ADDR_MASK4    32'h0000002b
`define NOC_NMU128__REG_ADDR_MASK4_SZ 32

`define NOC_NMU128__REG_ADDR_MASK5    32'h0000002c
`define NOC_NMU128__REG_ADDR_MASK5_SZ 32

`define NOC_NMU128__REG_ADDR_MASK6    32'h0000002d
`define NOC_NMU128__REG_ADDR_MASK6_SZ 32

`define NOC_NMU128__REG_ADDR_MASK7    32'h0000002e
`define NOC_NMU128__REG_ADDR_MASK7_SZ 32

`define NOC_NMU128__REG_ADDR_MASK8    32'h0000002f
`define NOC_NMU128__REG_ADDR_MASK8_SZ 32

`define NOC_NMU128__REG_ADDR_MASK9    32'h00000030
`define NOC_NMU128__REG_ADDR_MASK9_SZ 32

`define NOC_NMU128__REG_ADDR_REMAP    32'h00000031
`define NOC_NMU128__REG_ADDR_REMAP_SZ 16

`define NOC_NMU128__REG_ADDR_RPADDR0    32'h00000032
`define NOC_NMU128__REG_ADDR_RPADDR0_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR1    32'h00000033
`define NOC_NMU128__REG_ADDR_RPADDR1_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR10    32'h00000034
`define NOC_NMU128__REG_ADDR_RPADDR10_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR11    32'h00000035
`define NOC_NMU128__REG_ADDR_RPADDR11_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR12    32'h00000036
`define NOC_NMU128__REG_ADDR_RPADDR12_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR13    32'h00000037
`define NOC_NMU128__REG_ADDR_RPADDR13_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR14    32'h00000038
`define NOC_NMU128__REG_ADDR_RPADDR14_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR15    32'h00000039
`define NOC_NMU128__REG_ADDR_RPADDR15_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR2    32'h0000003a
`define NOC_NMU128__REG_ADDR_RPADDR2_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR3    32'h0000003b
`define NOC_NMU128__REG_ADDR_RPADDR3_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR4    32'h0000003c
`define NOC_NMU128__REG_ADDR_RPADDR4_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR5    32'h0000003d
`define NOC_NMU128__REG_ADDR_RPADDR5_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR6    32'h0000003e
`define NOC_NMU128__REG_ADDR_RPADDR6_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR7    32'h0000003f
`define NOC_NMU128__REG_ADDR_RPADDR7_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR8    32'h00000040
`define NOC_NMU128__REG_ADDR_RPADDR8_SZ 32

`define NOC_NMU128__REG_ADDR_RPADDR9    32'h00000041
`define NOC_NMU128__REG_ADDR_RPADDR9_SZ 32

`define NOC_NMU128__REG_ADR_MAP_CPM    32'h00000042
`define NOC_NMU128__REG_ADR_MAP_CPM_SZ 12

`define NOC_NMU128__REG_ADR_MAP_FPD_AFI_0    32'h00000043
`define NOC_NMU128__REG_ADR_MAP_FPD_AFI_0_SZ 12

`define NOC_NMU128__REG_ADR_MAP_FPD_AFI_1    32'h00000044
`define NOC_NMU128__REG_ADR_MAP_FPD_AFI_1_SZ 12

`define NOC_NMU128__REG_ADR_MAP_LPD_AFI_FS    32'h00000045
`define NOC_NMU128__REG_ADR_MAP_LPD_AFI_FS_SZ 12

`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_0    32'h00000046
`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_0_SZ 12

`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_1    32'h00000047
`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_1_SZ 12

`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_2    32'h00000048
`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_2_SZ 12

`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_3    32'h00000049
`define NOC_NMU128__REG_ADR_MAP_ME_ARRAY_3_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PCIE    32'h0000004a
`define NOC_NMU128__REG_ADR_MAP_PCIE_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PMC    32'h0000004b
`define NOC_NMU128__REG_ADR_MAP_PMC_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_0    32'h0000004c
`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_0_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_1    32'h0000004d
`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_1_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_2    32'h0000004e
`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_2_SZ 12

`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_3    32'h0000004f
`define NOC_NMU128__REG_ADR_MAP_PMC_ALIAS_3_SZ 12

`define NOC_NMU128__REG_ADR_MAP_QSPI    32'h00000050
`define NOC_NMU128__REG_ADR_MAP_QSPI_SZ 12

`define NOC_NMU128__REG_ADR_MAP_STM_GIC    32'h00000051
`define NOC_NMU128__REG_ADR_MAP_STM_GIC_SZ 12

`define NOC_NMU128__REG_ADR_MAP_XPDS    32'h00000052
`define NOC_NMU128__REG_ADR_MAP_XPDS_SZ 12

`define NOC_NMU128__REG_AXI_NON_MOD_DISABLE    32'h00000053
`define NOC_NMU128__REG_AXI_NON_MOD_DISABLE_SZ 1

`define NOC_NMU128__REG_AXI_PAR_CHK    32'h00000054
`define NOC_NMU128__REG_AXI_PAR_CHK_SZ 2

`define NOC_NMU128__REG_CHOPSIZE    32'h00000055
`define NOC_NMU128__REG_CHOPSIZE_SZ 4

`define NOC_NMU128__REG_DDR_ADR_MAP0    32'h00000056
`define NOC_NMU128__REG_DDR_ADR_MAP0_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP1    32'h00000057
`define NOC_NMU128__REG_DDR_ADR_MAP1_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP2    32'h00000058
`define NOC_NMU128__REG_DDR_ADR_MAP2_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP3    32'h00000059
`define NOC_NMU128__REG_DDR_ADR_MAP3_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP4    32'h0000005a
`define NOC_NMU128__REG_DDR_ADR_MAP4_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP5    32'h0000005b
`define NOC_NMU128__REG_DDR_ADR_MAP5_SZ 15

`define NOC_NMU128__REG_DDR_ADR_MAP6    32'h0000005c
`define NOC_NMU128__REG_DDR_ADR_MAP6_SZ 15

`define NOC_NMU128__REG_DDR_DST_MAP0    32'h0000005d
`define NOC_NMU128__REG_DDR_DST_MAP0_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP1    32'h0000005e
`define NOC_NMU128__REG_DDR_DST_MAP1_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP2    32'h0000005f
`define NOC_NMU128__REG_DDR_DST_MAP2_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP3    32'h00000060
`define NOC_NMU128__REG_DDR_DST_MAP3_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP4    32'h00000061
`define NOC_NMU128__REG_DDR_DST_MAP4_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP5    32'h00000062
`define NOC_NMU128__REG_DDR_DST_MAP5_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP6    32'h00000063
`define NOC_NMU128__REG_DDR_DST_MAP6_SZ 12

`define NOC_NMU128__REG_DDR_DST_MAP7    32'h00000064
`define NOC_NMU128__REG_DDR_DST_MAP7_SZ 12

`define NOC_NMU128__REG_DWIDTH    32'h00000065
`define NOC_NMU128__REG_DWIDTH_SZ 3

`define NOC_NMU128__REG_ECC_CHK_EN    32'h00000066
`define NOC_NMU128__REG_ECC_CHK_EN_SZ 1

`define NOC_NMU128__REG_HBM_MAP_T0_CH0    32'h00000067
`define NOC_NMU128__REG_HBM_MAP_T0_CH0_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH1    32'h00000068
`define NOC_NMU128__REG_HBM_MAP_T0_CH1_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH10    32'h00000069
`define NOC_NMU128__REG_HBM_MAP_T0_CH10_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH11    32'h0000006a
`define NOC_NMU128__REG_HBM_MAP_T0_CH11_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH12    32'h0000006b
`define NOC_NMU128__REG_HBM_MAP_T0_CH12_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH13    32'h0000006c
`define NOC_NMU128__REG_HBM_MAP_T0_CH13_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH14    32'h0000006d
`define NOC_NMU128__REG_HBM_MAP_T0_CH14_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH15    32'h0000006e
`define NOC_NMU128__REG_HBM_MAP_T0_CH15_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH2    32'h0000006f
`define NOC_NMU128__REG_HBM_MAP_T0_CH2_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH3    32'h00000070
`define NOC_NMU128__REG_HBM_MAP_T0_CH3_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH4    32'h00000071
`define NOC_NMU128__REG_HBM_MAP_T0_CH4_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH5    32'h00000072
`define NOC_NMU128__REG_HBM_MAP_T0_CH5_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH6    32'h00000073
`define NOC_NMU128__REG_HBM_MAP_T0_CH6_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH7    32'h00000074
`define NOC_NMU128__REG_HBM_MAP_T0_CH7_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH8    32'h00000075
`define NOC_NMU128__REG_HBM_MAP_T0_CH8_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T0_CH9    32'h00000076
`define NOC_NMU128__REG_HBM_MAP_T0_CH9_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH0    32'h00000077
`define NOC_NMU128__REG_HBM_MAP_T1_CH0_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH1    32'h00000078
`define NOC_NMU128__REG_HBM_MAP_T1_CH1_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH10    32'h00000079
`define NOC_NMU128__REG_HBM_MAP_T1_CH10_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH11    32'h0000007a
`define NOC_NMU128__REG_HBM_MAP_T1_CH11_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH12    32'h0000007b
`define NOC_NMU128__REG_HBM_MAP_T1_CH12_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH13    32'h0000007c
`define NOC_NMU128__REG_HBM_MAP_T1_CH13_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH14    32'h0000007d
`define NOC_NMU128__REG_HBM_MAP_T1_CH14_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH15    32'h0000007e
`define NOC_NMU128__REG_HBM_MAP_T1_CH15_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH2    32'h0000007f
`define NOC_NMU128__REG_HBM_MAP_T1_CH2_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH3    32'h00000080
`define NOC_NMU128__REG_HBM_MAP_T1_CH3_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH4    32'h00000081
`define NOC_NMU128__REG_HBM_MAP_T1_CH4_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH5    32'h00000082
`define NOC_NMU128__REG_HBM_MAP_T1_CH5_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH6    32'h00000083
`define NOC_NMU128__REG_HBM_MAP_T1_CH6_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH7    32'h00000084
`define NOC_NMU128__REG_HBM_MAP_T1_CH7_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH8    32'h00000085
`define NOC_NMU128__REG_HBM_MAP_T1_CH8_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T1_CH9    32'h00000086
`define NOC_NMU128__REG_HBM_MAP_T1_CH9_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH0    32'h00000087
`define NOC_NMU128__REG_HBM_MAP_T2_CH0_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH1    32'h00000088
`define NOC_NMU128__REG_HBM_MAP_T2_CH1_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH10    32'h00000089
`define NOC_NMU128__REG_HBM_MAP_T2_CH10_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH11    32'h0000008a
`define NOC_NMU128__REG_HBM_MAP_T2_CH11_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH12    32'h0000008b
`define NOC_NMU128__REG_HBM_MAP_T2_CH12_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH13    32'h0000008c
`define NOC_NMU128__REG_HBM_MAP_T2_CH13_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH14    32'h0000008d
`define NOC_NMU128__REG_HBM_MAP_T2_CH14_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH15    32'h0000008e
`define NOC_NMU128__REG_HBM_MAP_T2_CH15_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH2    32'h0000008f
`define NOC_NMU128__REG_HBM_MAP_T2_CH2_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH3    32'h00000090
`define NOC_NMU128__REG_HBM_MAP_T2_CH3_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH4    32'h00000091
`define NOC_NMU128__REG_HBM_MAP_T2_CH4_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH5    32'h00000092
`define NOC_NMU128__REG_HBM_MAP_T2_CH5_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH6    32'h00000093
`define NOC_NMU128__REG_HBM_MAP_T2_CH6_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH7    32'h00000094
`define NOC_NMU128__REG_HBM_MAP_T2_CH7_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH8    32'h00000095
`define NOC_NMU128__REG_HBM_MAP_T2_CH8_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T2_CH9    32'h00000096
`define NOC_NMU128__REG_HBM_MAP_T2_CH9_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH0    32'h00000097
`define NOC_NMU128__REG_HBM_MAP_T3_CH0_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH1    32'h00000098
`define NOC_NMU128__REG_HBM_MAP_T3_CH1_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH10    32'h00000099
`define NOC_NMU128__REG_HBM_MAP_T3_CH10_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH11    32'h0000009a
`define NOC_NMU128__REG_HBM_MAP_T3_CH11_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH12    32'h0000009b
`define NOC_NMU128__REG_HBM_MAP_T3_CH12_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH13    32'h0000009c
`define NOC_NMU128__REG_HBM_MAP_T3_CH13_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH14    32'h0000009d
`define NOC_NMU128__REG_HBM_MAP_T3_CH14_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH15    32'h0000009e
`define NOC_NMU128__REG_HBM_MAP_T3_CH15_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH2    32'h0000009f
`define NOC_NMU128__REG_HBM_MAP_T3_CH2_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH3    32'h000000a0
`define NOC_NMU128__REG_HBM_MAP_T3_CH3_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH4    32'h000000a1
`define NOC_NMU128__REG_HBM_MAP_T3_CH4_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH5    32'h000000a2
`define NOC_NMU128__REG_HBM_MAP_T3_CH5_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH6    32'h000000a3
`define NOC_NMU128__REG_HBM_MAP_T3_CH6_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH7    32'h000000a4
`define NOC_NMU128__REG_HBM_MAP_T3_CH7_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH8    32'h000000a5
`define NOC_NMU128__REG_HBM_MAP_T3_CH8_SZ 12

`define NOC_NMU128__REG_HBM_MAP_T3_CH9    32'h000000a6
`define NOC_NMU128__REG_HBM_MAP_T3_CH9_SZ 12

`define NOC_NMU128__REG_MODE_SELECT    32'h000000a7
`define NOC_NMU128__REG_MODE_SELECT_SZ 16

`define NOC_NMU128__REG_OUTSTANDING_RD_TXN    32'h000000a8
`define NOC_NMU128__REG_OUTSTANDING_RD_TXN_SZ 7

`define NOC_NMU128__REG_OUTSTANDING_WR_TXN    32'h000000a9
`define NOC_NMU128__REG_OUTSTANDING_WR_TXN_SZ 7

`define NOC_NMU128__REG_PRIORITY    32'h000000aa
`define NOC_NMU128__REG_PRIORITY_SZ 2

`define NOC_NMU128__REG_RD_AXPROT_SEL    32'h000000ab
`define NOC_NMU128__REG_RD_AXPROT_SEL_SZ 6

`define NOC_NMU128__REG_RD_RATE_CREDIT_DROP    32'h000000ac
`define NOC_NMU128__REG_RD_RATE_CREDIT_DROP_SZ 10

`define NOC_NMU128__REG_RD_RATE_CREDIT_LIMIT    32'h000000ad
`define NOC_NMU128__REG_RD_RATE_CREDIT_LIMIT_SZ 13

`define NOC_NMU128__REG_RD_VCA_TOKEN0    32'h000000ae
`define NOC_NMU128__REG_RD_VCA_TOKEN0_SZ 8

`define NOC_NMU128__REG_RPOISON_TO_SLVERR    32'h000000af
`define NOC_NMU128__REG_RPOISON_TO_SLVERR_SZ 1

`define NOC_NMU128__REG_RROB_RAM_SETTING    32'h000000b0
`define NOC_NMU128__REG_RROB_RAM_SETTING_SZ 9

`define NOC_NMU128__REG_SMID_SEL    32'h000000b1
`define NOC_NMU128__REG_SMID_SEL_SZ 20

`define NOC_NMU128__REG_SRC    32'h000000b2
`define NOC_NMU128__REG_SRC_SZ 12

`define NOC_NMU128__REG_TBASE_AXI_TIMEOUT    32'h000000b3
`define NOC_NMU128__REG_TBASE_AXI_TIMEOUT_SZ 4

`define NOC_NMU128__REG_TBASE_MODE_RLIMIT_RD    32'h000000b4
`define NOC_NMU128__REG_TBASE_MODE_RLIMIT_RD_SZ 3

`define NOC_NMU128__REG_TBASE_MODE_RLIMIT_WR    32'h000000b5
`define NOC_NMU128__REG_TBASE_MODE_RLIMIT_WR_SZ 3

`define NOC_NMU128__REG_TBASE_TRK_TIMEOUT    32'h000000b6
`define NOC_NMU128__REG_TBASE_TRK_TIMEOUT_SZ 4

`define NOC_NMU128__REG_VC_MAP    32'h000000b7
`define NOC_NMU128__REG_VC_MAP_SZ 12

`define NOC_NMU128__REG_WBUF_LAUNCH_SIZE    32'h000000b8
`define NOC_NMU128__REG_WBUF_LAUNCH_SIZE_SZ 6

`define NOC_NMU128__REG_WBUF_RAM_SETTING    32'h000000b9
`define NOC_NMU128__REG_WBUF_RAM_SETTING_SZ 9

`define NOC_NMU128__REG_WR_AXPROT_SEL    32'h000000ba
`define NOC_NMU128__REG_WR_AXPROT_SEL_SZ 6

`define NOC_NMU128__REG_WR_RATE_CREDIT_DROP    32'h000000bb
`define NOC_NMU128__REG_WR_RATE_CREDIT_DROP_SZ 10

`define NOC_NMU128__REG_WR_RATE_CREDIT_LIMIT    32'h000000bc
`define NOC_NMU128__REG_WR_RATE_CREDIT_LIMIT_SZ 13

`define NOC_NMU128__REG_WR_VCA_TOKEN0    32'h000000bd
`define NOC_NMU128__REG_WR_VCA_TOKEN0_SZ 8

`endif  // B_NOC_NMU128_DEFINES_VH