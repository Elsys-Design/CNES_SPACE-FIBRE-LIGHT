// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IOBUFDS_INTERMDISABLE_ODDR_DEFINES_VH
`else
`define B_IOBUFDS_INTERMDISABLE_ODDR_DEFINES_VH

// Look-up table parameters
//

`define IOBUFDS_INTERMDISABLE_ODDR_ADDR_N  4
`define IOBUFDS_INTERMDISABLE_ODDR_ADDR_SZ 32
`define IOBUFDS_INTERMDISABLE_ODDR_DATA_SZ 56

// Attribute addresses
//

`define IOBUFDS_INTERMDISABLE_ODDR__DIFF_TERM    32'h00000000
`define IOBUFDS_INTERMDISABLE_ODDR__DIFF_TERM_SZ 40

`define IOBUFDS_INTERMDISABLE_ODDR__DQS_BIAS    32'h00000001
`define IOBUFDS_INTERMDISABLE_ODDR__DQS_BIAS_SZ 40

`define IOBUFDS_INTERMDISABLE_ODDR__IOSTANDARD    32'h00000002
`define IOBUFDS_INTERMDISABLE_ODDR__IOSTANDARD_SZ 56

`define IOBUFDS_INTERMDISABLE_ODDR__USE_IBUFDISABLE    32'h00000003
`define IOBUFDS_INTERMDISABLE_ODDR__USE_IBUFDISABLE_SZ 40

`endif  // B_IOBUFDS_INTERMDISABLE_ODDR_DEFINES_VH