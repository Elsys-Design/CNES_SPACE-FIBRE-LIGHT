// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC_NPS6_DEFINES_VH
`else
`define B_NOC_NPS6_DEFINES_VH

// Look-up table parameters
//

`define NOC_NPS6_ADDR_N  559
`define NOC_NPS6_ADDR_SZ 32
`define NOC_NPS6_DATA_SZ 32

// Attribute addresses
//

`define NOC_NPS6__REG_CLOCK_MUX    32'h00000000
`define NOC_NPS6__REG_CLOCK_MUX_SZ 32

`define NOC_NPS6__REG_HIGH_ID0_P0    32'h00000001
`define NOC_NPS6__REG_HIGH_ID0_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID0_P1    32'h00000002
`define NOC_NPS6__REG_HIGH_ID0_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID0_P2    32'h00000003
`define NOC_NPS6__REG_HIGH_ID0_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID0_P3    32'h00000004
`define NOC_NPS6__REG_HIGH_ID0_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID0_P4    32'h00000005
`define NOC_NPS6__REG_HIGH_ID0_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID0_P5    32'h00000006
`define NOC_NPS6__REG_HIGH_ID0_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID10_P0    32'h00000007
`define NOC_NPS6__REG_HIGH_ID10_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID10_P1    32'h00000008
`define NOC_NPS6__REG_HIGH_ID10_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID10_P2    32'h00000009
`define NOC_NPS6__REG_HIGH_ID10_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID10_P3    32'h0000000a
`define NOC_NPS6__REG_HIGH_ID10_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID10_P4    32'h0000000b
`define NOC_NPS6__REG_HIGH_ID10_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID10_P5    32'h0000000c
`define NOC_NPS6__REG_HIGH_ID10_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID11_P0    32'h0000000d
`define NOC_NPS6__REG_HIGH_ID11_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID11_P1    32'h0000000e
`define NOC_NPS6__REG_HIGH_ID11_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID11_P2    32'h0000000f
`define NOC_NPS6__REG_HIGH_ID11_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID11_P3    32'h00000010
`define NOC_NPS6__REG_HIGH_ID11_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID11_P4    32'h00000011
`define NOC_NPS6__REG_HIGH_ID11_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID11_P5    32'h00000012
`define NOC_NPS6__REG_HIGH_ID11_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID12_P0    32'h00000013
`define NOC_NPS6__REG_HIGH_ID12_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID12_P1    32'h00000014
`define NOC_NPS6__REG_HIGH_ID12_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID12_P2    32'h00000015
`define NOC_NPS6__REG_HIGH_ID12_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID12_P3    32'h00000016
`define NOC_NPS6__REG_HIGH_ID12_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID12_P4    32'h00000017
`define NOC_NPS6__REG_HIGH_ID12_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID12_P5    32'h00000018
`define NOC_NPS6__REG_HIGH_ID12_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID13_P0    32'h00000019
`define NOC_NPS6__REG_HIGH_ID13_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID13_P1    32'h0000001a
`define NOC_NPS6__REG_HIGH_ID13_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID13_P2    32'h0000001b
`define NOC_NPS6__REG_HIGH_ID13_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID13_P3    32'h0000001c
`define NOC_NPS6__REG_HIGH_ID13_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID13_P4    32'h0000001d
`define NOC_NPS6__REG_HIGH_ID13_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID13_P5    32'h0000001e
`define NOC_NPS6__REG_HIGH_ID13_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID14_P0    32'h0000001f
`define NOC_NPS6__REG_HIGH_ID14_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID14_P1    32'h00000020
`define NOC_NPS6__REG_HIGH_ID14_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID14_P2    32'h00000021
`define NOC_NPS6__REG_HIGH_ID14_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID14_P3    32'h00000022
`define NOC_NPS6__REG_HIGH_ID14_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID14_P4    32'h00000023
`define NOC_NPS6__REG_HIGH_ID14_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID14_P5    32'h00000024
`define NOC_NPS6__REG_HIGH_ID14_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID15_P0    32'h00000025
`define NOC_NPS6__REG_HIGH_ID15_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID15_P1    32'h00000026
`define NOC_NPS6__REG_HIGH_ID15_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID15_P2    32'h00000027
`define NOC_NPS6__REG_HIGH_ID15_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID15_P3    32'h00000028
`define NOC_NPS6__REG_HIGH_ID15_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID15_P4    32'h00000029
`define NOC_NPS6__REG_HIGH_ID15_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID15_P5    32'h0000002a
`define NOC_NPS6__REG_HIGH_ID15_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID16_P0    32'h0000002b
`define NOC_NPS6__REG_HIGH_ID16_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID16_P1    32'h0000002c
`define NOC_NPS6__REG_HIGH_ID16_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID16_P2    32'h0000002d
`define NOC_NPS6__REG_HIGH_ID16_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID16_P3    32'h0000002e
`define NOC_NPS6__REG_HIGH_ID16_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID16_P4    32'h0000002f
`define NOC_NPS6__REG_HIGH_ID16_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID16_P5    32'h00000030
`define NOC_NPS6__REG_HIGH_ID16_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID17_P0    32'h00000031
`define NOC_NPS6__REG_HIGH_ID17_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID17_P1    32'h00000032
`define NOC_NPS6__REG_HIGH_ID17_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID17_P2    32'h00000033
`define NOC_NPS6__REG_HIGH_ID17_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID17_P3    32'h00000034
`define NOC_NPS6__REG_HIGH_ID17_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID17_P4    32'h00000035
`define NOC_NPS6__REG_HIGH_ID17_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID17_P5    32'h00000036
`define NOC_NPS6__REG_HIGH_ID17_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID18_P0    32'h00000037
`define NOC_NPS6__REG_HIGH_ID18_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID18_P1    32'h00000038
`define NOC_NPS6__REG_HIGH_ID18_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID18_P2    32'h00000039
`define NOC_NPS6__REG_HIGH_ID18_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID18_P3    32'h0000003a
`define NOC_NPS6__REG_HIGH_ID18_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID18_P4    32'h0000003b
`define NOC_NPS6__REG_HIGH_ID18_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID18_P5    32'h0000003c
`define NOC_NPS6__REG_HIGH_ID18_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID19_P0    32'h0000003d
`define NOC_NPS6__REG_HIGH_ID19_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID19_P1    32'h0000003e
`define NOC_NPS6__REG_HIGH_ID19_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID19_P2    32'h0000003f
`define NOC_NPS6__REG_HIGH_ID19_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID19_P3    32'h00000040
`define NOC_NPS6__REG_HIGH_ID19_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID19_P4    32'h00000041
`define NOC_NPS6__REG_HIGH_ID19_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID19_P5    32'h00000042
`define NOC_NPS6__REG_HIGH_ID19_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID1_P0    32'h00000043
`define NOC_NPS6__REG_HIGH_ID1_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID1_P1    32'h00000044
`define NOC_NPS6__REG_HIGH_ID1_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID1_P2    32'h00000045
`define NOC_NPS6__REG_HIGH_ID1_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID1_P3    32'h00000046
`define NOC_NPS6__REG_HIGH_ID1_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID1_P4    32'h00000047
`define NOC_NPS6__REG_HIGH_ID1_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID1_P5    32'h00000048
`define NOC_NPS6__REG_HIGH_ID1_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID20_P0    32'h00000049
`define NOC_NPS6__REG_HIGH_ID20_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID20_P1    32'h0000004a
`define NOC_NPS6__REG_HIGH_ID20_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID20_P2    32'h0000004b
`define NOC_NPS6__REG_HIGH_ID20_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID20_P3    32'h0000004c
`define NOC_NPS6__REG_HIGH_ID20_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID20_P4    32'h0000004d
`define NOC_NPS6__REG_HIGH_ID20_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID20_P5    32'h0000004e
`define NOC_NPS6__REG_HIGH_ID20_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID21_P0    32'h0000004f
`define NOC_NPS6__REG_HIGH_ID21_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID21_P1    32'h00000050
`define NOC_NPS6__REG_HIGH_ID21_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID21_P2    32'h00000051
`define NOC_NPS6__REG_HIGH_ID21_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID21_P3    32'h00000052
`define NOC_NPS6__REG_HIGH_ID21_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID21_P4    32'h00000053
`define NOC_NPS6__REG_HIGH_ID21_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID21_P5    32'h00000054
`define NOC_NPS6__REG_HIGH_ID21_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID22_P0    32'h00000055
`define NOC_NPS6__REG_HIGH_ID22_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID22_P1    32'h00000056
`define NOC_NPS6__REG_HIGH_ID22_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID22_P2    32'h00000057
`define NOC_NPS6__REG_HIGH_ID22_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID22_P3    32'h00000058
`define NOC_NPS6__REG_HIGH_ID22_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID22_P4    32'h00000059
`define NOC_NPS6__REG_HIGH_ID22_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID22_P5    32'h0000005a
`define NOC_NPS6__REG_HIGH_ID22_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID23_P0    32'h0000005b
`define NOC_NPS6__REG_HIGH_ID23_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID23_P1    32'h0000005c
`define NOC_NPS6__REG_HIGH_ID23_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID23_P2    32'h0000005d
`define NOC_NPS6__REG_HIGH_ID23_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID23_P3    32'h0000005e
`define NOC_NPS6__REG_HIGH_ID23_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID23_P4    32'h0000005f
`define NOC_NPS6__REG_HIGH_ID23_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID23_P5    32'h00000060
`define NOC_NPS6__REG_HIGH_ID23_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID24_P0    32'h00000061
`define NOC_NPS6__REG_HIGH_ID24_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID24_P1    32'h00000062
`define NOC_NPS6__REG_HIGH_ID24_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID24_P2    32'h00000063
`define NOC_NPS6__REG_HIGH_ID24_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID24_P3    32'h00000064
`define NOC_NPS6__REG_HIGH_ID24_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID24_P4    32'h00000065
`define NOC_NPS6__REG_HIGH_ID24_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID24_P5    32'h00000066
`define NOC_NPS6__REG_HIGH_ID24_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID25_P0    32'h00000067
`define NOC_NPS6__REG_HIGH_ID25_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID25_P1    32'h00000068
`define NOC_NPS6__REG_HIGH_ID25_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID25_P2    32'h00000069
`define NOC_NPS6__REG_HIGH_ID25_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID25_P3    32'h0000006a
`define NOC_NPS6__REG_HIGH_ID25_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID25_P4    32'h0000006b
`define NOC_NPS6__REG_HIGH_ID25_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID25_P5    32'h0000006c
`define NOC_NPS6__REG_HIGH_ID25_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID26_P0    32'h0000006d
`define NOC_NPS6__REG_HIGH_ID26_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID26_P1    32'h0000006e
`define NOC_NPS6__REG_HIGH_ID26_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID26_P2    32'h0000006f
`define NOC_NPS6__REG_HIGH_ID26_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID26_P3    32'h00000070
`define NOC_NPS6__REG_HIGH_ID26_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID26_P4    32'h00000071
`define NOC_NPS6__REG_HIGH_ID26_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID26_P5    32'h00000072
`define NOC_NPS6__REG_HIGH_ID26_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID27_P0    32'h00000073
`define NOC_NPS6__REG_HIGH_ID27_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID27_P1    32'h00000074
`define NOC_NPS6__REG_HIGH_ID27_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID27_P2    32'h00000075
`define NOC_NPS6__REG_HIGH_ID27_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID27_P3    32'h00000076
`define NOC_NPS6__REG_HIGH_ID27_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID27_P4    32'h00000077
`define NOC_NPS6__REG_HIGH_ID27_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID27_P5    32'h00000078
`define NOC_NPS6__REG_HIGH_ID27_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID28_P0    32'h00000079
`define NOC_NPS6__REG_HIGH_ID28_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID28_P1    32'h0000007a
`define NOC_NPS6__REG_HIGH_ID28_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID28_P2    32'h0000007b
`define NOC_NPS6__REG_HIGH_ID28_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID28_P3    32'h0000007c
`define NOC_NPS6__REG_HIGH_ID28_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID28_P4    32'h0000007d
`define NOC_NPS6__REG_HIGH_ID28_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID28_P5    32'h0000007e
`define NOC_NPS6__REG_HIGH_ID28_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID29_P0    32'h0000007f
`define NOC_NPS6__REG_HIGH_ID29_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID29_P1    32'h00000080
`define NOC_NPS6__REG_HIGH_ID29_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID29_P2    32'h00000081
`define NOC_NPS6__REG_HIGH_ID29_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID29_P3    32'h00000082
`define NOC_NPS6__REG_HIGH_ID29_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID29_P4    32'h00000083
`define NOC_NPS6__REG_HIGH_ID29_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID29_P5    32'h00000084
`define NOC_NPS6__REG_HIGH_ID29_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID2_P0    32'h00000085
`define NOC_NPS6__REG_HIGH_ID2_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID2_P1    32'h00000086
`define NOC_NPS6__REG_HIGH_ID2_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID2_P2    32'h00000087
`define NOC_NPS6__REG_HIGH_ID2_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID2_P3    32'h00000088
`define NOC_NPS6__REG_HIGH_ID2_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID2_P4    32'h00000089
`define NOC_NPS6__REG_HIGH_ID2_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID2_P5    32'h0000008a
`define NOC_NPS6__REG_HIGH_ID2_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID30_P0    32'h0000008b
`define NOC_NPS6__REG_HIGH_ID30_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID30_P1    32'h0000008c
`define NOC_NPS6__REG_HIGH_ID30_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID30_P2    32'h0000008d
`define NOC_NPS6__REG_HIGH_ID30_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID30_P3    32'h0000008e
`define NOC_NPS6__REG_HIGH_ID30_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID30_P4    32'h0000008f
`define NOC_NPS6__REG_HIGH_ID30_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID30_P5    32'h00000090
`define NOC_NPS6__REG_HIGH_ID30_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID31_P0    32'h00000091
`define NOC_NPS6__REG_HIGH_ID31_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID31_P1    32'h00000092
`define NOC_NPS6__REG_HIGH_ID31_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID31_P2    32'h00000093
`define NOC_NPS6__REG_HIGH_ID31_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID31_P3    32'h00000094
`define NOC_NPS6__REG_HIGH_ID31_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID31_P4    32'h00000095
`define NOC_NPS6__REG_HIGH_ID31_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID31_P5    32'h00000096
`define NOC_NPS6__REG_HIGH_ID31_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID32_P0    32'h00000097
`define NOC_NPS6__REG_HIGH_ID32_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID32_P1    32'h00000098
`define NOC_NPS6__REG_HIGH_ID32_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID32_P2    32'h00000099
`define NOC_NPS6__REG_HIGH_ID32_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID32_P3    32'h0000009a
`define NOC_NPS6__REG_HIGH_ID32_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID32_P4    32'h0000009b
`define NOC_NPS6__REG_HIGH_ID32_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID32_P5    32'h0000009c
`define NOC_NPS6__REG_HIGH_ID32_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID33_P0    32'h0000009d
`define NOC_NPS6__REG_HIGH_ID33_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID33_P1    32'h0000009e
`define NOC_NPS6__REG_HIGH_ID33_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID33_P2    32'h0000009f
`define NOC_NPS6__REG_HIGH_ID33_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID33_P3    32'h000000a0
`define NOC_NPS6__REG_HIGH_ID33_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID33_P4    32'h000000a1
`define NOC_NPS6__REG_HIGH_ID33_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID33_P5    32'h000000a2
`define NOC_NPS6__REG_HIGH_ID33_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID34_P0    32'h000000a3
`define NOC_NPS6__REG_HIGH_ID34_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID34_P1    32'h000000a4
`define NOC_NPS6__REG_HIGH_ID34_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID34_P2    32'h000000a5
`define NOC_NPS6__REG_HIGH_ID34_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID34_P3    32'h000000a6
`define NOC_NPS6__REG_HIGH_ID34_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID34_P4    32'h000000a7
`define NOC_NPS6__REG_HIGH_ID34_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID34_P5    32'h000000a8
`define NOC_NPS6__REG_HIGH_ID34_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID35_P0    32'h000000a9
`define NOC_NPS6__REG_HIGH_ID35_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID35_P1    32'h000000aa
`define NOC_NPS6__REG_HIGH_ID35_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID35_P2    32'h000000ab
`define NOC_NPS6__REG_HIGH_ID35_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID35_P3    32'h000000ac
`define NOC_NPS6__REG_HIGH_ID35_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID35_P4    32'h000000ad
`define NOC_NPS6__REG_HIGH_ID35_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID35_P5    32'h000000ae
`define NOC_NPS6__REG_HIGH_ID35_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID36_P0    32'h000000af
`define NOC_NPS6__REG_HIGH_ID36_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID36_P1    32'h000000b0
`define NOC_NPS6__REG_HIGH_ID36_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID36_P2    32'h000000b1
`define NOC_NPS6__REG_HIGH_ID36_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID36_P3    32'h000000b2
`define NOC_NPS6__REG_HIGH_ID36_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID36_P4    32'h000000b3
`define NOC_NPS6__REG_HIGH_ID36_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID36_P5    32'h000000b4
`define NOC_NPS6__REG_HIGH_ID36_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID37_P0    32'h000000b5
`define NOC_NPS6__REG_HIGH_ID37_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID37_P1    32'h000000b6
`define NOC_NPS6__REG_HIGH_ID37_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID37_P2    32'h000000b7
`define NOC_NPS6__REG_HIGH_ID37_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID37_P3    32'h000000b8
`define NOC_NPS6__REG_HIGH_ID37_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID37_P4    32'h000000b9
`define NOC_NPS6__REG_HIGH_ID37_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID37_P5    32'h000000ba
`define NOC_NPS6__REG_HIGH_ID37_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID38_P0    32'h000000bb
`define NOC_NPS6__REG_HIGH_ID38_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID38_P1    32'h000000bc
`define NOC_NPS6__REG_HIGH_ID38_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID38_P2    32'h000000bd
`define NOC_NPS6__REG_HIGH_ID38_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID38_P3    32'h000000be
`define NOC_NPS6__REG_HIGH_ID38_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID38_P4    32'h000000bf
`define NOC_NPS6__REG_HIGH_ID38_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID38_P5    32'h000000c0
`define NOC_NPS6__REG_HIGH_ID38_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID39_P0    32'h000000c1
`define NOC_NPS6__REG_HIGH_ID39_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID39_P1    32'h000000c2
`define NOC_NPS6__REG_HIGH_ID39_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID39_P2    32'h000000c3
`define NOC_NPS6__REG_HIGH_ID39_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID39_P3    32'h000000c4
`define NOC_NPS6__REG_HIGH_ID39_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID39_P4    32'h000000c5
`define NOC_NPS6__REG_HIGH_ID39_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID39_P5    32'h000000c6
`define NOC_NPS6__REG_HIGH_ID39_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID3_P0    32'h000000c7
`define NOC_NPS6__REG_HIGH_ID3_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID3_P1    32'h000000c8
`define NOC_NPS6__REG_HIGH_ID3_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID3_P2    32'h000000c9
`define NOC_NPS6__REG_HIGH_ID3_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID3_P3    32'h000000ca
`define NOC_NPS6__REG_HIGH_ID3_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID3_P4    32'h000000cb
`define NOC_NPS6__REG_HIGH_ID3_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID3_P5    32'h000000cc
`define NOC_NPS6__REG_HIGH_ID3_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID40_P0    32'h000000cd
`define NOC_NPS6__REG_HIGH_ID40_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID40_P1    32'h000000ce
`define NOC_NPS6__REG_HIGH_ID40_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID40_P2    32'h000000cf
`define NOC_NPS6__REG_HIGH_ID40_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID40_P3    32'h000000d0
`define NOC_NPS6__REG_HIGH_ID40_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID40_P4    32'h000000d1
`define NOC_NPS6__REG_HIGH_ID40_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID40_P5    32'h000000d2
`define NOC_NPS6__REG_HIGH_ID40_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID41_P0    32'h000000d3
`define NOC_NPS6__REG_HIGH_ID41_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID41_P1    32'h000000d4
`define NOC_NPS6__REG_HIGH_ID41_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID41_P2    32'h000000d5
`define NOC_NPS6__REG_HIGH_ID41_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID41_P3    32'h000000d6
`define NOC_NPS6__REG_HIGH_ID41_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID41_P4    32'h000000d7
`define NOC_NPS6__REG_HIGH_ID41_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID41_P5    32'h000000d8
`define NOC_NPS6__REG_HIGH_ID41_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID42_P0    32'h000000d9
`define NOC_NPS6__REG_HIGH_ID42_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID42_P1    32'h000000da
`define NOC_NPS6__REG_HIGH_ID42_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID42_P2    32'h000000db
`define NOC_NPS6__REG_HIGH_ID42_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID42_P3    32'h000000dc
`define NOC_NPS6__REG_HIGH_ID42_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID42_P4    32'h000000dd
`define NOC_NPS6__REG_HIGH_ID42_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID42_P5    32'h000000de
`define NOC_NPS6__REG_HIGH_ID42_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID43_P0    32'h000000df
`define NOC_NPS6__REG_HIGH_ID43_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID43_P1    32'h000000e0
`define NOC_NPS6__REG_HIGH_ID43_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID43_P2    32'h000000e1
`define NOC_NPS6__REG_HIGH_ID43_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID43_P3    32'h000000e2
`define NOC_NPS6__REG_HIGH_ID43_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID43_P4    32'h000000e3
`define NOC_NPS6__REG_HIGH_ID43_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID43_P5    32'h000000e4
`define NOC_NPS6__REG_HIGH_ID43_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID44_P0    32'h000000e5
`define NOC_NPS6__REG_HIGH_ID44_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID44_P1    32'h000000e6
`define NOC_NPS6__REG_HIGH_ID44_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID44_P2    32'h000000e7
`define NOC_NPS6__REG_HIGH_ID44_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID44_P3    32'h000000e8
`define NOC_NPS6__REG_HIGH_ID44_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID44_P4    32'h000000e9
`define NOC_NPS6__REG_HIGH_ID44_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID44_P5    32'h000000ea
`define NOC_NPS6__REG_HIGH_ID44_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID45_P0    32'h000000eb
`define NOC_NPS6__REG_HIGH_ID45_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID45_P1    32'h000000ec
`define NOC_NPS6__REG_HIGH_ID45_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID45_P2    32'h000000ed
`define NOC_NPS6__REG_HIGH_ID45_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID45_P3    32'h000000ee
`define NOC_NPS6__REG_HIGH_ID45_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID45_P4    32'h000000ef
`define NOC_NPS6__REG_HIGH_ID45_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID45_P5    32'h000000f0
`define NOC_NPS6__REG_HIGH_ID45_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID46_P0    32'h000000f1
`define NOC_NPS6__REG_HIGH_ID46_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID46_P1    32'h000000f2
`define NOC_NPS6__REG_HIGH_ID46_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID46_P2    32'h000000f3
`define NOC_NPS6__REG_HIGH_ID46_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID46_P3    32'h000000f4
`define NOC_NPS6__REG_HIGH_ID46_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID46_P4    32'h000000f5
`define NOC_NPS6__REG_HIGH_ID46_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID46_P5    32'h000000f6
`define NOC_NPS6__REG_HIGH_ID46_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID47_P0    32'h000000f7
`define NOC_NPS6__REG_HIGH_ID47_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID47_P1    32'h000000f8
`define NOC_NPS6__REG_HIGH_ID47_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID47_P2    32'h000000f9
`define NOC_NPS6__REG_HIGH_ID47_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID47_P3    32'h000000fa
`define NOC_NPS6__REG_HIGH_ID47_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID47_P4    32'h000000fb
`define NOC_NPS6__REG_HIGH_ID47_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID47_P5    32'h000000fc
`define NOC_NPS6__REG_HIGH_ID47_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID48_P0    32'h000000fd
`define NOC_NPS6__REG_HIGH_ID48_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID48_P1    32'h000000fe
`define NOC_NPS6__REG_HIGH_ID48_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID48_P2    32'h000000ff
`define NOC_NPS6__REG_HIGH_ID48_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID48_P3    32'h00000100
`define NOC_NPS6__REG_HIGH_ID48_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID48_P4    32'h00000101
`define NOC_NPS6__REG_HIGH_ID48_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID48_P5    32'h00000102
`define NOC_NPS6__REG_HIGH_ID48_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID49_P0    32'h00000103
`define NOC_NPS6__REG_HIGH_ID49_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID49_P1    32'h00000104
`define NOC_NPS6__REG_HIGH_ID49_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID49_P2    32'h00000105
`define NOC_NPS6__REG_HIGH_ID49_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID49_P3    32'h00000106
`define NOC_NPS6__REG_HIGH_ID49_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID49_P4    32'h00000107
`define NOC_NPS6__REG_HIGH_ID49_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID49_P5    32'h00000108
`define NOC_NPS6__REG_HIGH_ID49_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID4_P0    32'h00000109
`define NOC_NPS6__REG_HIGH_ID4_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID4_P1    32'h0000010a
`define NOC_NPS6__REG_HIGH_ID4_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID4_P2    32'h0000010b
`define NOC_NPS6__REG_HIGH_ID4_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID4_P3    32'h0000010c
`define NOC_NPS6__REG_HIGH_ID4_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID4_P4    32'h0000010d
`define NOC_NPS6__REG_HIGH_ID4_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID4_P5    32'h0000010e
`define NOC_NPS6__REG_HIGH_ID4_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID50_P0    32'h0000010f
`define NOC_NPS6__REG_HIGH_ID50_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID50_P1    32'h00000110
`define NOC_NPS6__REG_HIGH_ID50_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID50_P2    32'h00000111
`define NOC_NPS6__REG_HIGH_ID50_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID50_P3    32'h00000112
`define NOC_NPS6__REG_HIGH_ID50_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID50_P4    32'h00000113
`define NOC_NPS6__REG_HIGH_ID50_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID50_P5    32'h00000114
`define NOC_NPS6__REG_HIGH_ID50_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID51_P0    32'h00000115
`define NOC_NPS6__REG_HIGH_ID51_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID51_P1    32'h00000116
`define NOC_NPS6__REG_HIGH_ID51_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID51_P2    32'h00000117
`define NOC_NPS6__REG_HIGH_ID51_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID51_P3    32'h00000118
`define NOC_NPS6__REG_HIGH_ID51_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID51_P4    32'h00000119
`define NOC_NPS6__REG_HIGH_ID51_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID51_P5    32'h0000011a
`define NOC_NPS6__REG_HIGH_ID51_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID52_P0    32'h0000011b
`define NOC_NPS6__REG_HIGH_ID52_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID52_P1    32'h0000011c
`define NOC_NPS6__REG_HIGH_ID52_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID52_P2    32'h0000011d
`define NOC_NPS6__REG_HIGH_ID52_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID52_P3    32'h0000011e
`define NOC_NPS6__REG_HIGH_ID52_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID52_P4    32'h0000011f
`define NOC_NPS6__REG_HIGH_ID52_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID52_P5    32'h00000120
`define NOC_NPS6__REG_HIGH_ID52_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID53_P0    32'h00000121
`define NOC_NPS6__REG_HIGH_ID53_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID53_P1    32'h00000122
`define NOC_NPS6__REG_HIGH_ID53_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID53_P2    32'h00000123
`define NOC_NPS6__REG_HIGH_ID53_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID53_P3    32'h00000124
`define NOC_NPS6__REG_HIGH_ID53_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID53_P4    32'h00000125
`define NOC_NPS6__REG_HIGH_ID53_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID53_P5    32'h00000126
`define NOC_NPS6__REG_HIGH_ID53_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID54_P0    32'h00000127
`define NOC_NPS6__REG_HIGH_ID54_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID54_P1    32'h00000128
`define NOC_NPS6__REG_HIGH_ID54_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID54_P2    32'h00000129
`define NOC_NPS6__REG_HIGH_ID54_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID54_P3    32'h0000012a
`define NOC_NPS6__REG_HIGH_ID54_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID54_P4    32'h0000012b
`define NOC_NPS6__REG_HIGH_ID54_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID54_P5    32'h0000012c
`define NOC_NPS6__REG_HIGH_ID54_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID55_P0    32'h0000012d
`define NOC_NPS6__REG_HIGH_ID55_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID55_P1    32'h0000012e
`define NOC_NPS6__REG_HIGH_ID55_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID55_P2    32'h0000012f
`define NOC_NPS6__REG_HIGH_ID55_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID55_P3    32'h00000130
`define NOC_NPS6__REG_HIGH_ID55_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID55_P4    32'h00000131
`define NOC_NPS6__REG_HIGH_ID55_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID55_P5    32'h00000132
`define NOC_NPS6__REG_HIGH_ID55_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID56_P0    32'h00000133
`define NOC_NPS6__REG_HIGH_ID56_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID56_P1    32'h00000134
`define NOC_NPS6__REG_HIGH_ID56_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID56_P2    32'h00000135
`define NOC_NPS6__REG_HIGH_ID56_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID56_P3    32'h00000136
`define NOC_NPS6__REG_HIGH_ID56_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID56_P4    32'h00000137
`define NOC_NPS6__REG_HIGH_ID56_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID56_P5    32'h00000138
`define NOC_NPS6__REG_HIGH_ID56_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID57_P0    32'h00000139
`define NOC_NPS6__REG_HIGH_ID57_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID57_P1    32'h0000013a
`define NOC_NPS6__REG_HIGH_ID57_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID57_P2    32'h0000013b
`define NOC_NPS6__REG_HIGH_ID57_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID57_P3    32'h0000013c
`define NOC_NPS6__REG_HIGH_ID57_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID57_P4    32'h0000013d
`define NOC_NPS6__REG_HIGH_ID57_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID57_P5    32'h0000013e
`define NOC_NPS6__REG_HIGH_ID57_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID58_P0    32'h0000013f
`define NOC_NPS6__REG_HIGH_ID58_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID58_P1    32'h00000140
`define NOC_NPS6__REG_HIGH_ID58_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID58_P2    32'h00000141
`define NOC_NPS6__REG_HIGH_ID58_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID58_P3    32'h00000142
`define NOC_NPS6__REG_HIGH_ID58_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID58_P4    32'h00000143
`define NOC_NPS6__REG_HIGH_ID58_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID58_P5    32'h00000144
`define NOC_NPS6__REG_HIGH_ID58_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID59_P0    32'h00000145
`define NOC_NPS6__REG_HIGH_ID59_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID59_P1    32'h00000146
`define NOC_NPS6__REG_HIGH_ID59_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID59_P2    32'h00000147
`define NOC_NPS6__REG_HIGH_ID59_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID59_P3    32'h00000148
`define NOC_NPS6__REG_HIGH_ID59_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID59_P4    32'h00000149
`define NOC_NPS6__REG_HIGH_ID59_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID59_P5    32'h0000014a
`define NOC_NPS6__REG_HIGH_ID59_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID5_P0    32'h0000014b
`define NOC_NPS6__REG_HIGH_ID5_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID5_P1    32'h0000014c
`define NOC_NPS6__REG_HIGH_ID5_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID5_P2    32'h0000014d
`define NOC_NPS6__REG_HIGH_ID5_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID5_P3    32'h0000014e
`define NOC_NPS6__REG_HIGH_ID5_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID5_P4    32'h0000014f
`define NOC_NPS6__REG_HIGH_ID5_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID5_P5    32'h00000150
`define NOC_NPS6__REG_HIGH_ID5_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID60_P0    32'h00000151
`define NOC_NPS6__REG_HIGH_ID60_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID60_P1    32'h00000152
`define NOC_NPS6__REG_HIGH_ID60_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID60_P2    32'h00000153
`define NOC_NPS6__REG_HIGH_ID60_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID60_P3    32'h00000154
`define NOC_NPS6__REG_HIGH_ID60_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID60_P4    32'h00000155
`define NOC_NPS6__REG_HIGH_ID60_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID60_P5    32'h00000156
`define NOC_NPS6__REG_HIGH_ID60_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID61_P0    32'h00000157
`define NOC_NPS6__REG_HIGH_ID61_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID61_P1    32'h00000158
`define NOC_NPS6__REG_HIGH_ID61_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID61_P2    32'h00000159
`define NOC_NPS6__REG_HIGH_ID61_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID61_P3    32'h0000015a
`define NOC_NPS6__REG_HIGH_ID61_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID61_P4    32'h0000015b
`define NOC_NPS6__REG_HIGH_ID61_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID61_P5    32'h0000015c
`define NOC_NPS6__REG_HIGH_ID61_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID62_P0    32'h0000015d
`define NOC_NPS6__REG_HIGH_ID62_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID62_P1    32'h0000015e
`define NOC_NPS6__REG_HIGH_ID62_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID62_P2    32'h0000015f
`define NOC_NPS6__REG_HIGH_ID62_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID62_P3    32'h00000160
`define NOC_NPS6__REG_HIGH_ID62_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID62_P4    32'h00000161
`define NOC_NPS6__REG_HIGH_ID62_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID62_P5    32'h00000162
`define NOC_NPS6__REG_HIGH_ID62_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID63_P0    32'h00000163
`define NOC_NPS6__REG_HIGH_ID63_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID63_P1    32'h00000164
`define NOC_NPS6__REG_HIGH_ID63_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID63_P2    32'h00000165
`define NOC_NPS6__REG_HIGH_ID63_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID63_P3    32'h00000166
`define NOC_NPS6__REG_HIGH_ID63_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID63_P4    32'h00000167
`define NOC_NPS6__REG_HIGH_ID63_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID63_P5    32'h00000168
`define NOC_NPS6__REG_HIGH_ID63_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID6_P0    32'h00000169
`define NOC_NPS6__REG_HIGH_ID6_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID6_P1    32'h0000016a
`define NOC_NPS6__REG_HIGH_ID6_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID6_P2    32'h0000016b
`define NOC_NPS6__REG_HIGH_ID6_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID6_P3    32'h0000016c
`define NOC_NPS6__REG_HIGH_ID6_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID6_P4    32'h0000016d
`define NOC_NPS6__REG_HIGH_ID6_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID6_P5    32'h0000016e
`define NOC_NPS6__REG_HIGH_ID6_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID7_P0    32'h0000016f
`define NOC_NPS6__REG_HIGH_ID7_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID7_P1    32'h00000170
`define NOC_NPS6__REG_HIGH_ID7_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID7_P2    32'h00000171
`define NOC_NPS6__REG_HIGH_ID7_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID7_P3    32'h00000172
`define NOC_NPS6__REG_HIGH_ID7_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID7_P4    32'h00000173
`define NOC_NPS6__REG_HIGH_ID7_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID7_P5    32'h00000174
`define NOC_NPS6__REG_HIGH_ID7_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID8_P0    32'h00000175
`define NOC_NPS6__REG_HIGH_ID8_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID8_P1    32'h00000176
`define NOC_NPS6__REG_HIGH_ID8_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID8_P2    32'h00000177
`define NOC_NPS6__REG_HIGH_ID8_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID8_P3    32'h00000178
`define NOC_NPS6__REG_HIGH_ID8_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID8_P4    32'h00000179
`define NOC_NPS6__REG_HIGH_ID8_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID8_P5    32'h0000017a
`define NOC_NPS6__REG_HIGH_ID8_P5_SZ 31

`define NOC_NPS6__REG_HIGH_ID9_P0    32'h0000017b
`define NOC_NPS6__REG_HIGH_ID9_P0_SZ 31

`define NOC_NPS6__REG_HIGH_ID9_P1    32'h0000017c
`define NOC_NPS6__REG_HIGH_ID9_P1_SZ 23

`define NOC_NPS6__REG_HIGH_ID9_P2    32'h0000017d
`define NOC_NPS6__REG_HIGH_ID9_P2_SZ 23

`define NOC_NPS6__REG_HIGH_ID9_P3    32'h0000017e
`define NOC_NPS6__REG_HIGH_ID9_P3_SZ 31

`define NOC_NPS6__REG_HIGH_ID9_P4    32'h0000017f
`define NOC_NPS6__REG_HIGH_ID9_P4_SZ 31

`define NOC_NPS6__REG_HIGH_ID9_P5    32'h00000180
`define NOC_NPS6__REG_HIGH_ID9_P5_SZ 31

`define NOC_NPS6__REG_ID    32'h00000181
`define NOC_NPS6__REG_ID_SZ 10

`define NOC_NPS6__REG_LOW_ID0_P0    32'h00000182
`define NOC_NPS6__REG_LOW_ID0_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID0_P1    32'h00000183
`define NOC_NPS6__REG_LOW_ID0_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID0_P2    32'h00000184
`define NOC_NPS6__REG_LOW_ID0_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID0_P3    32'h00000185
`define NOC_NPS6__REG_LOW_ID0_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID0_P4    32'h00000186
`define NOC_NPS6__REG_LOW_ID0_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID0_P5    32'h00000187
`define NOC_NPS6__REG_LOW_ID0_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID10_P0    32'h00000188
`define NOC_NPS6__REG_LOW_ID10_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID10_P1    32'h00000189
`define NOC_NPS6__REG_LOW_ID10_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID10_P2    32'h0000018a
`define NOC_NPS6__REG_LOW_ID10_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID10_P3    32'h0000018b
`define NOC_NPS6__REG_LOW_ID10_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID10_P4    32'h0000018c
`define NOC_NPS6__REG_LOW_ID10_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID10_P5    32'h0000018d
`define NOC_NPS6__REG_LOW_ID10_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID11_P0    32'h0000018e
`define NOC_NPS6__REG_LOW_ID11_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID11_P1    32'h0000018f
`define NOC_NPS6__REG_LOW_ID11_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID11_P2    32'h00000190
`define NOC_NPS6__REG_LOW_ID11_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID11_P3    32'h00000191
`define NOC_NPS6__REG_LOW_ID11_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID11_P4    32'h00000192
`define NOC_NPS6__REG_LOW_ID11_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID11_P5    32'h00000193
`define NOC_NPS6__REG_LOW_ID11_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID12_P0    32'h00000194
`define NOC_NPS6__REG_LOW_ID12_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID12_P1    32'h00000195
`define NOC_NPS6__REG_LOW_ID12_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID12_P2    32'h00000196
`define NOC_NPS6__REG_LOW_ID12_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID12_P3    32'h00000197
`define NOC_NPS6__REG_LOW_ID12_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID12_P4    32'h00000198
`define NOC_NPS6__REG_LOW_ID12_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID12_P5    32'h00000199
`define NOC_NPS6__REG_LOW_ID12_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID13_P0    32'h0000019a
`define NOC_NPS6__REG_LOW_ID13_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID13_P1    32'h0000019b
`define NOC_NPS6__REG_LOW_ID13_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID13_P2    32'h0000019c
`define NOC_NPS6__REG_LOW_ID13_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID13_P3    32'h0000019d
`define NOC_NPS6__REG_LOW_ID13_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID13_P4    32'h0000019e
`define NOC_NPS6__REG_LOW_ID13_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID13_P5    32'h0000019f
`define NOC_NPS6__REG_LOW_ID13_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID14_P0    32'h000001a0
`define NOC_NPS6__REG_LOW_ID14_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID14_P1    32'h000001a1
`define NOC_NPS6__REG_LOW_ID14_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID14_P2    32'h000001a2
`define NOC_NPS6__REG_LOW_ID14_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID14_P3    32'h000001a3
`define NOC_NPS6__REG_LOW_ID14_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID14_P4    32'h000001a4
`define NOC_NPS6__REG_LOW_ID14_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID14_P5    32'h000001a5
`define NOC_NPS6__REG_LOW_ID14_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID15_P0    32'h000001a6
`define NOC_NPS6__REG_LOW_ID15_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID15_P1    32'h000001a7
`define NOC_NPS6__REG_LOW_ID15_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID15_P2    32'h000001a8
`define NOC_NPS6__REG_LOW_ID15_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID15_P3    32'h000001a9
`define NOC_NPS6__REG_LOW_ID15_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID15_P4    32'h000001aa
`define NOC_NPS6__REG_LOW_ID15_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID15_P5    32'h000001ab
`define NOC_NPS6__REG_LOW_ID15_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID1_P0    32'h000001ac
`define NOC_NPS6__REG_LOW_ID1_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID1_P1    32'h000001ad
`define NOC_NPS6__REG_LOW_ID1_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID1_P2    32'h000001ae
`define NOC_NPS6__REG_LOW_ID1_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID1_P3    32'h000001af
`define NOC_NPS6__REG_LOW_ID1_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID1_P4    32'h000001b0
`define NOC_NPS6__REG_LOW_ID1_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID1_P5    32'h000001b1
`define NOC_NPS6__REG_LOW_ID1_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID2_P0    32'h000001b2
`define NOC_NPS6__REG_LOW_ID2_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID2_P1    32'h000001b3
`define NOC_NPS6__REG_LOW_ID2_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID2_P2    32'h000001b4
`define NOC_NPS6__REG_LOW_ID2_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID2_P3    32'h000001b5
`define NOC_NPS6__REG_LOW_ID2_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID2_P4    32'h000001b6
`define NOC_NPS6__REG_LOW_ID2_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID2_P5    32'h000001b7
`define NOC_NPS6__REG_LOW_ID2_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID3_P0    32'h000001b8
`define NOC_NPS6__REG_LOW_ID3_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID3_P1    32'h000001b9
`define NOC_NPS6__REG_LOW_ID3_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID3_P2    32'h000001ba
`define NOC_NPS6__REG_LOW_ID3_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID3_P3    32'h000001bb
`define NOC_NPS6__REG_LOW_ID3_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID3_P4    32'h000001bc
`define NOC_NPS6__REG_LOW_ID3_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID3_P5    32'h000001bd
`define NOC_NPS6__REG_LOW_ID3_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID4_P0    32'h000001be
`define NOC_NPS6__REG_LOW_ID4_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID4_P1    32'h000001bf
`define NOC_NPS6__REG_LOW_ID4_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID4_P2    32'h000001c0
`define NOC_NPS6__REG_LOW_ID4_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID4_P3    32'h000001c1
`define NOC_NPS6__REG_LOW_ID4_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID4_P4    32'h000001c2
`define NOC_NPS6__REG_LOW_ID4_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID4_P5    32'h000001c3
`define NOC_NPS6__REG_LOW_ID4_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID5_P0    32'h000001c4
`define NOC_NPS6__REG_LOW_ID5_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID5_P1    32'h000001c5
`define NOC_NPS6__REG_LOW_ID5_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID5_P2    32'h000001c6
`define NOC_NPS6__REG_LOW_ID5_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID5_P3    32'h000001c7
`define NOC_NPS6__REG_LOW_ID5_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID5_P4    32'h000001c8
`define NOC_NPS6__REG_LOW_ID5_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID5_P5    32'h000001c9
`define NOC_NPS6__REG_LOW_ID5_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID6_P0    32'h000001ca
`define NOC_NPS6__REG_LOW_ID6_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID6_P1    32'h000001cb
`define NOC_NPS6__REG_LOW_ID6_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID6_P2    32'h000001cc
`define NOC_NPS6__REG_LOW_ID6_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID6_P3    32'h000001cd
`define NOC_NPS6__REG_LOW_ID6_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID6_P4    32'h000001ce
`define NOC_NPS6__REG_LOW_ID6_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID6_P5    32'h000001cf
`define NOC_NPS6__REG_LOW_ID6_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID7_P0    32'h000001d0
`define NOC_NPS6__REG_LOW_ID7_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID7_P1    32'h000001d1
`define NOC_NPS6__REG_LOW_ID7_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID7_P2    32'h000001d2
`define NOC_NPS6__REG_LOW_ID7_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID7_P3    32'h000001d3
`define NOC_NPS6__REG_LOW_ID7_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID7_P4    32'h000001d4
`define NOC_NPS6__REG_LOW_ID7_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID7_P5    32'h000001d5
`define NOC_NPS6__REG_LOW_ID7_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID8_P0    32'h000001d6
`define NOC_NPS6__REG_LOW_ID8_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID8_P1    32'h000001d7
`define NOC_NPS6__REG_LOW_ID8_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID8_P2    32'h000001d8
`define NOC_NPS6__REG_LOW_ID8_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID8_P3    32'h000001d9
`define NOC_NPS6__REG_LOW_ID8_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID8_P4    32'h000001da
`define NOC_NPS6__REG_LOW_ID8_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID8_P5    32'h000001db
`define NOC_NPS6__REG_LOW_ID8_P5_SZ 31

`define NOC_NPS6__REG_LOW_ID9_P0    32'h000001dc
`define NOC_NPS6__REG_LOW_ID9_P0_SZ 31

`define NOC_NPS6__REG_LOW_ID9_P1    32'h000001dd
`define NOC_NPS6__REG_LOW_ID9_P1_SZ 23

`define NOC_NPS6__REG_LOW_ID9_P2    32'h000001de
`define NOC_NPS6__REG_LOW_ID9_P2_SZ 23

`define NOC_NPS6__REG_LOW_ID9_P3    32'h000001df
`define NOC_NPS6__REG_LOW_ID9_P3_SZ 31

`define NOC_NPS6__REG_LOW_ID9_P4    32'h000001e0
`define NOC_NPS6__REG_LOW_ID9_P4_SZ 31

`define NOC_NPS6__REG_LOW_ID9_P5    32'h000001e1
`define NOC_NPS6__REG_LOW_ID9_P5_SZ 31

`define NOC_NPS6__REG_MID_ID0_P0    32'h000001e2
`define NOC_NPS6__REG_MID_ID0_P0_SZ 31

`define NOC_NPS6__REG_MID_ID0_P1    32'h000001e3
`define NOC_NPS6__REG_MID_ID0_P1_SZ 23

`define NOC_NPS6__REG_MID_ID0_P2    32'h000001e4
`define NOC_NPS6__REG_MID_ID0_P2_SZ 23

`define NOC_NPS6__REG_MID_ID0_P3    32'h000001e5
`define NOC_NPS6__REG_MID_ID0_P3_SZ 31

`define NOC_NPS6__REG_MID_ID0_P4    32'h000001e6
`define NOC_NPS6__REG_MID_ID0_P4_SZ 31

`define NOC_NPS6__REG_MID_ID0_P5    32'h000001e7
`define NOC_NPS6__REG_MID_ID0_P5_SZ 31

`define NOC_NPS6__REG_MID_ID1_P0    32'h000001e8
`define NOC_NPS6__REG_MID_ID1_P0_SZ 31

`define NOC_NPS6__REG_MID_ID1_P1    32'h000001e9
`define NOC_NPS6__REG_MID_ID1_P1_SZ 23

`define NOC_NPS6__REG_MID_ID1_P2    32'h000001ea
`define NOC_NPS6__REG_MID_ID1_P2_SZ 23

`define NOC_NPS6__REG_MID_ID1_P3    32'h000001eb
`define NOC_NPS6__REG_MID_ID1_P3_SZ 31

`define NOC_NPS6__REG_MID_ID1_P4    32'h000001ec
`define NOC_NPS6__REG_MID_ID1_P4_SZ 31

`define NOC_NPS6__REG_MID_ID1_P5    32'h000001ed
`define NOC_NPS6__REG_MID_ID1_P5_SZ 31

`define NOC_NPS6__REG_MID_ID2_P0    32'h000001ee
`define NOC_NPS6__REG_MID_ID2_P0_SZ 31

`define NOC_NPS6__REG_MID_ID2_P1    32'h000001ef
`define NOC_NPS6__REG_MID_ID2_P1_SZ 23

`define NOC_NPS6__REG_MID_ID2_P2    32'h000001f0
`define NOC_NPS6__REG_MID_ID2_P2_SZ 23

`define NOC_NPS6__REG_MID_ID2_P3    32'h000001f1
`define NOC_NPS6__REG_MID_ID2_P3_SZ 31

`define NOC_NPS6__REG_MID_ID2_P4    32'h000001f2
`define NOC_NPS6__REG_MID_ID2_P4_SZ 31

`define NOC_NPS6__REG_MID_ID2_P5    32'h000001f3
`define NOC_NPS6__REG_MID_ID2_P5_SZ 31

`define NOC_NPS6__REG_MID_ID3_P0    32'h000001f4
`define NOC_NPS6__REG_MID_ID3_P0_SZ 31

`define NOC_NPS6__REG_MID_ID3_P1    32'h000001f5
`define NOC_NPS6__REG_MID_ID3_P1_SZ 23

`define NOC_NPS6__REG_MID_ID3_P2    32'h000001f6
`define NOC_NPS6__REG_MID_ID3_P2_SZ 23

`define NOC_NPS6__REG_MID_ID3_P3    32'h000001f7
`define NOC_NPS6__REG_MID_ID3_P3_SZ 31

`define NOC_NPS6__REG_MID_ID3_P4    32'h000001f8
`define NOC_NPS6__REG_MID_ID3_P4_SZ 31

`define NOC_NPS6__REG_MID_ID3_P5    32'h000001f9
`define NOC_NPS6__REG_MID_ID3_P5_SZ 31

`define NOC_NPS6__REG_NOC_CTL    32'h000001fa
`define NOC_NPS6__REG_NOC_CTL_SZ 16

`define NOC_NPS6__REG_P00_P1_0_VCA_TOKEN    32'h000001fb
`define NOC_NPS6__REG_P00_P1_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P00_P1_1_VCA_TOKEN    32'h000001fc
`define NOC_NPS6__REG_P00_P1_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P01_P2_0_VCA_TOKEN    32'h000001fd
`define NOC_NPS6__REG_P01_P2_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P01_P2_1_VCA_TOKEN    32'h000001fe
`define NOC_NPS6__REG_P01_P2_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P02_P3_0_VCA_TOKEN    32'h000001ff
`define NOC_NPS6__REG_P02_P3_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P02_P3_1_VCA_TOKEN    32'h00000200
`define NOC_NPS6__REG_P02_P3_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P03_P4_0_VCA_TOKEN    32'h00000201
`define NOC_NPS6__REG_P03_P4_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P03_P4_1_VCA_TOKEN    32'h00000202
`define NOC_NPS6__REG_P03_P4_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P04_P5_0_VCA_TOKEN    32'h00000203
`define NOC_NPS6__REG_P04_P5_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P04_P5_1_VCA_TOKEN    32'h00000204
`define NOC_NPS6__REG_P04_P5_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P10_P3_0_VCA_TOKEN    32'h00000205
`define NOC_NPS6__REG_P10_P3_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P10_P3_1_VCA_TOKEN    32'h00000206
`define NOC_NPS6__REG_P10_P3_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P11_P4_0_VCA_TOKEN    32'h00000207
`define NOC_NPS6__REG_P11_P4_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P11_P4_1_VCA_TOKEN    32'h00000208
`define NOC_NPS6__REG_P11_P4_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P12_P5_0_VCA_TOKEN    32'h00000209
`define NOC_NPS6__REG_P12_P5_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P12_P5_1_VCA_TOKEN    32'h0000020a
`define NOC_NPS6__REG_P12_P5_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P13_P0_0_VCA_TOKEN    32'h0000020b
`define NOC_NPS6__REG_P13_P0_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P13_P0_1_VCA_TOKEN    32'h0000020c
`define NOC_NPS6__REG_P13_P0_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P20_P4_0_VCA_TOKEN    32'h0000020d
`define NOC_NPS6__REG_P20_P4_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P20_P4_1_VCA_TOKEN    32'h0000020e
`define NOC_NPS6__REG_P20_P4_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P21_P5_0_VCA_TOKEN    32'h0000020f
`define NOC_NPS6__REG_P21_P5_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P21_P5_1_VCA_TOKEN    32'h00000210
`define NOC_NPS6__REG_P21_P5_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P22_P0_0_VCA_TOKEN    32'h00000211
`define NOC_NPS6__REG_P22_P0_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P22_P0_1_VCA_TOKEN    32'h00000212
`define NOC_NPS6__REG_P22_P0_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P23_P3_0_VCA_TOKEN    32'h00000213
`define NOC_NPS6__REG_P23_P3_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P23_P3_1_VCA_TOKEN    32'h00000214
`define NOC_NPS6__REG_P23_P3_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P30_P5_0_VCA_TOKEN    32'h00000215
`define NOC_NPS6__REG_P30_P5_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P30_P5_1_VCA_TOKEN    32'h00000216
`define NOC_NPS6__REG_P30_P5_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P31_P0_0_VCA_TOKEN    32'h00000217
`define NOC_NPS6__REG_P31_P0_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P31_P0_1_VCA_TOKEN    32'h00000218
`define NOC_NPS6__REG_P31_P0_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P32_P1_0_VCA_TOKEN    32'h00000219
`define NOC_NPS6__REG_P32_P1_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P32_P1_1_VCA_TOKEN    32'h0000021a
`define NOC_NPS6__REG_P32_P1_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P33_P2_0_VCA_TOKEN    32'h0000021b
`define NOC_NPS6__REG_P33_P2_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P33_P2_1_VCA_TOKEN    32'h0000021c
`define NOC_NPS6__REG_P33_P2_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P34_P4_0_VCA_TOKEN    32'h0000021d
`define NOC_NPS6__REG_P34_P4_0_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P34_P4_1_VCA_TOKEN    32'h0000021e
`define NOC_NPS6__REG_P34_P4_1_VCA_TOKEN_SZ 32

`define NOC_NPS6__REG_P40_P0_0_VCA_TOKEN    32'h0000021f
`define NOC_NPS6__REG_P40_P0_0_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P40_P0_1_VCA_TOKEN    32'h00000220
`define NOC_NPS6__REG_P40_P0_1_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P41_P1_0_VCA_TOKEN    32'h00000221
`define NOC_NPS6__REG_P41_P1_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P41_P1_1_VCA_TOKEN    32'h00000222
`define NOC_NPS6__REG_P41_P1_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P42_P2_0_VCA_TOKEN    32'h00000223
`define NOC_NPS6__REG_P42_P2_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P42_P2_1_VCA_TOKEN    32'h00000224
`define NOC_NPS6__REG_P42_P2_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P43_P3_0_VCA_TOKEN    32'h00000225
`define NOC_NPS6__REG_P43_P3_0_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P43_P3_1_VCA_TOKEN    32'h00000226
`define NOC_NPS6__REG_P43_P3_1_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P50_P1_0_VCA_TOKEN    32'h00000227
`define NOC_NPS6__REG_P50_P1_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P50_P1_1_VCA_TOKEN    32'h00000228
`define NOC_NPS6__REG_P50_P1_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P51_P2_0_VCA_TOKEN    32'h00000229
`define NOC_NPS6__REG_P51_P2_0_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P51_P2_1_VCA_TOKEN    32'h0000022a
`define NOC_NPS6__REG_P51_P2_1_VCA_TOKEN_SZ 16

`define NOC_NPS6__REG_P52_P3_0_VCA_TOKEN    32'h0000022b
`define NOC_NPS6__REG_P52_P3_0_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P52_P3_1_VCA_TOKEN    32'h0000022c
`define NOC_NPS6__REG_P52_P3_1_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P53_P0_0_VCA_TOKEN    32'h0000022d
`define NOC_NPS6__REG_P53_P0_0_VCA_TOKEN_SZ 24

`define NOC_NPS6__REG_P53_P0_1_VCA_TOKEN    32'h0000022e
`define NOC_NPS6__REG_P53_P0_1_VCA_TOKEN_SZ 24

`endif  // B_NOC_NPS6_DEFINES_VH