`include "B_BUFGCE_DIV_defines.vh"

reg [`BUFGCE_DIV_DATA_SZ-1:0] ATTR [0:`BUFGCE_DIV_ADDR_N-1];
reg [`BUFGCE_DIV__BUFGCE_DIVIDE_SZ-1:0] BUFGCE_DIVIDE_REG = BUFGCE_DIVIDE;
reg [`BUFGCE_DIV__CE_TYPE_SZ:1] CE_TYPE_REG = CE_TYPE;
reg [`BUFGCE_DIV__HARDSYNC_CLR_SZ:1] HARDSYNC_CLR_REG = HARDSYNC_CLR;
reg IS_CE_INVERTED_REG = IS_CE_INVERTED;
reg IS_CLR_INVERTED_REG = IS_CLR_INVERTED;
reg IS_I_INVERTED_REG = IS_I_INVERTED;
reg [`BUFGCE_DIV__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`BUFGCE_DIV__STARTUP_SYNC_SZ:1] STARTUP_SYNC_REG = STARTUP_SYNC;

initial begin
  ATTR[`BUFGCE_DIV__BUFGCE_DIVIDE] = BUFGCE_DIVIDE;
  ATTR[`BUFGCE_DIV__CE_TYPE] = CE_TYPE;
  ATTR[`BUFGCE_DIV__HARDSYNC_CLR] = HARDSYNC_CLR;
  ATTR[`BUFGCE_DIV__IS_CE_INVERTED] = IS_CE_INVERTED;
  ATTR[`BUFGCE_DIV__IS_CLR_INVERTED] = IS_CLR_INVERTED;
  ATTR[`BUFGCE_DIV__IS_I_INVERTED] = IS_I_INVERTED;
  ATTR[`BUFGCE_DIV__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`BUFGCE_DIV__STARTUP_SYNC] = STARTUP_SYNC;
end

always @(trig_attr) begin
  BUFGCE_DIVIDE_REG = ATTR[`BUFGCE_DIV__BUFGCE_DIVIDE];
  CE_TYPE_REG = ATTR[`BUFGCE_DIV__CE_TYPE];
  HARDSYNC_CLR_REG = ATTR[`BUFGCE_DIV__HARDSYNC_CLR];
  IS_CE_INVERTED_REG = ATTR[`BUFGCE_DIV__IS_CE_INVERTED];
  IS_CLR_INVERTED_REG = ATTR[`BUFGCE_DIV__IS_CLR_INVERTED];
  IS_I_INVERTED_REG = ATTR[`BUFGCE_DIV__IS_I_INVERTED];
  SIM_DEVICE_REG = ATTR[`BUFGCE_DIV__SIM_DEVICE];
  STARTUP_SYNC_REG = ATTR[`BUFGCE_DIV__STARTUP_SYNC];
end

// procedures to override, read attribute values

task write_attr;
  input  [`BUFGCE_DIV_ADDR_SZ-1:0] addr;
  input  [`BUFGCE_DIV_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`BUFGCE_DIV_DATA_SZ-1:0] read_attr;
  input  [`BUFGCE_DIV_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
