// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_ALU_DEFINES_VH
`else
`define B_DSP_ALU_DEFINES_VH

// Look-up table parameters
//

`define DSP_ALU_ADDR_N  16
`define DSP_ALU_ADDR_SZ 32
`define DSP_ALU_DATA_SZ 88

// Attribute addresses
//

`define DSP_ALU__ALUMODEREG    32'h00000000
`define DSP_ALU__ALUMODEREG_SZ 32

`define DSP_ALU__CARRYINREG    32'h00000001
`define DSP_ALU__CARRYINREG_SZ 32

`define DSP_ALU__CARRYINSELREG    32'h00000002
`define DSP_ALU__CARRYINSELREG_SZ 32

`define DSP_ALU__IS_ALUMODE_INVERTED    32'h00000003
`define DSP_ALU__IS_ALUMODE_INVERTED_SZ 4

`define DSP_ALU__IS_CARRYIN_INVERTED    32'h00000004
`define DSP_ALU__IS_CARRYIN_INVERTED_SZ 1

`define DSP_ALU__IS_CLK_INVERTED    32'h00000005
`define DSP_ALU__IS_CLK_INVERTED_SZ 1

`define DSP_ALU__IS_OPMODE_INVERTED    32'h00000006
`define DSP_ALU__IS_OPMODE_INVERTED_SZ 9

`define DSP_ALU__IS_RSTALLCARRYIN_INVERTED    32'h00000007
`define DSP_ALU__IS_RSTALLCARRYIN_INVERTED_SZ 1

`define DSP_ALU__IS_RSTALUMODE_INVERTED    32'h00000008
`define DSP_ALU__IS_RSTALUMODE_INVERTED_SZ 1

`define DSP_ALU__IS_RSTCTRL_INVERTED    32'h00000009
`define DSP_ALU__IS_RSTCTRL_INVERTED_SZ 1

`define DSP_ALU__MREG    32'h0000000a
`define DSP_ALU__MREG_SZ 32

`define DSP_ALU__OPMODEREG    32'h0000000b
`define DSP_ALU__OPMODEREG_SZ 32

`define DSP_ALU__RND    32'h0000000c
`define DSP_ALU__RND_SZ 48

`define DSP_ALU__USE_SIMD    32'h0000000d
`define DSP_ALU__USE_SIMD_SZ 48

`define DSP_ALU__USE_WIDEXOR    32'h0000000e
`define DSP_ALU__USE_WIDEXOR_SZ 40

`define DSP_ALU__XORSIMD    32'h0000000f
`define DSP_ALU__XORSIMD_SZ 88

`endif  // B_DSP_ALU_DEFINES_VH