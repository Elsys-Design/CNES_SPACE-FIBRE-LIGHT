// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP48E1_DEFINES_VH
`else
`define B_DSP48E1_DEFINES_VH

// Look-up table parameters
//

`define DSP48E1_ADDR_N  30
`define DSP48E1_ADDR_SZ 32
`define DSP48E1_DATA_SZ 120

// Attribute addresses
//

`define DSP48E1__ACASCREG    32'h00000000
`define DSP48E1__ACASCREG_SZ 32

`define DSP48E1__ADREG    32'h00000001
`define DSP48E1__ADREG_SZ 32

`define DSP48E1__ALUMODEREG    32'h00000002
`define DSP48E1__ALUMODEREG_SZ 32

`define DSP48E1__AREG    32'h00000003
`define DSP48E1__AREG_SZ 32

`define DSP48E1__AUTORESET_PATDET    32'h00000004
`define DSP48E1__AUTORESET_PATDET_SZ 120

`define DSP48E1__A_INPUT    32'h00000005
`define DSP48E1__A_INPUT_SZ 56

`define DSP48E1__BCASCREG    32'h00000006
`define DSP48E1__BCASCREG_SZ 32

`define DSP48E1__BREG    32'h00000007
`define DSP48E1__BREG_SZ 32

`define DSP48E1__B_INPUT    32'h00000008
`define DSP48E1__B_INPUT_SZ 56

`define DSP48E1__CARRYINREG    32'h00000009
`define DSP48E1__CARRYINREG_SZ 32

`define DSP48E1__CARRYINSELREG    32'h0000000a
`define DSP48E1__CARRYINSELREG_SZ 32

`define DSP48E1__CREG    32'h0000000b
`define DSP48E1__CREG_SZ 32

`define DSP48E1__DREG    32'h0000000c
`define DSP48E1__DREG_SZ 32

`define DSP48E1__INMODEREG    32'h0000000d
`define DSP48E1__INMODEREG_SZ 32

`define DSP48E1__IS_ALUMODE_INVERTED    32'h0000000e
`define DSP48E1__IS_ALUMODE_INVERTED_SZ 4

`define DSP48E1__IS_CARRYIN_INVERTED    32'h0000000f
`define DSP48E1__IS_CARRYIN_INVERTED_SZ 1

`define DSP48E1__IS_CLK_INVERTED    32'h00000010
`define DSP48E1__IS_CLK_INVERTED_SZ 1

`define DSP48E1__IS_INMODE_INVERTED    32'h00000011
`define DSP48E1__IS_INMODE_INVERTED_SZ 5

`define DSP48E1__IS_OPMODE_INVERTED    32'h00000012
`define DSP48E1__IS_OPMODE_INVERTED_SZ 7

`define DSP48E1__MASK    32'h00000013
`define DSP48E1__MASK_SZ 48

`define DSP48E1__MREG    32'h00000014
`define DSP48E1__MREG_SZ 32

`define DSP48E1__OPMODEREG    32'h00000015
`define DSP48E1__OPMODEREG_SZ 32

`define DSP48E1__PATTERN    32'h00000016
`define DSP48E1__PATTERN_SZ 48

`define DSP48E1__PREG    32'h00000017
`define DSP48E1__PREG_SZ 32

`define DSP48E1__SEL_MASK    32'h00000018
`define DSP48E1__SEL_MASK_SZ 112

`define DSP48E1__SEL_PATTERN    32'h00000019
`define DSP48E1__SEL_PATTERN_SZ 56

`define DSP48E1__USE_DPORT    32'h0000001a
`define DSP48E1__USE_DPORT_SZ 40

`define DSP48E1__USE_MULT    32'h0000001b
`define DSP48E1__USE_MULT_SZ 64

`define DSP48E1__USE_PATTERN_DETECT    32'h0000001c
`define DSP48E1__USE_PATTERN_DETECT_SZ 72

`define DSP48E1__USE_SIMD    32'h0000001d
`define DSP48E1__USE_SIMD_SZ 48

`endif  // B_DSP48E1_DEFINES_VH