--------------------------------------------------------------------------
-- COMPANY       : ELSYS Design
--------------------------------------------------------------------------
-- TITLE         : lane_configurator.vhd
-- PROJECT       : SPACE FIBRE LIGHT
--------------------------------------------------------------------------
-- AUTHOR        : Yvan DAURIAC
-- CREATED       : 31/08/2024
--------------------------------------------------------------------------
-- DESCRIPTION   : Model able to communicate with IP PHY/LANE MIB blocks
--------------------------------------------------------------------------
-- History       : V1.0: Creation of the file
--------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_model.all;
------------------------------------------------------------------------------------------------------------------
--                                                      ENTITY                                                  --
------------------------------------------------------------------------------------------------------------------
entity LANE_CONFIGURATOR is
    generic(
       G_ADDR_WIDTH : positive := C_AXI_ADDR_WIDTH;                              -- Generic for AXI address width
       G_DATA_WIDTH : positive := C_AXI_DATA_WIDTH                               -- Generic for AXI data width
    );
    port(
   -- Clock and reset
   ------------------
   CLK                   : in std_logic;                                         -- Clock signal
   RST_N                 : in std_logic;                                         -- Reset active low signal
   CLK_TX                : in  std_logic;                                        -- Clock generated by manufacturer IP
   RST_TXCLK_N           : in  std_logic;                                        -- Reset clock generated by manufacturer IP
   -- AXI4 Lite slave interface
   ---------------------------------------
       -- Write Address channel (AW)
   S_AXI_AWADDR          : in std_logic_vector(G_ADDR_WIDTH-1 downto 0);         -- Write address from master to slave
   S_AXI_AWVALID         : in std_logic;                                         -- Master asserts when write address is valid
   S_AXI_AWREADY         : out std_logic;                                        -- Slave ready to accept write address
       -- Write Data channel (W)
   S_AXI_WDATA           : in std_logic_vector(G_DATA_WIDTH-1 downto 0);         -- Write data from master
   S_AXI_WSTRB           : in std_logic_vector(3 downto 0);                      -- Write strobe, indicates active byte lanes
   S_AXI_WVALID          : in std_logic;                                         -- Master asserts when write data is valid
   S_AXI_WREADY          : out std_logic;                                        -- Slave ready to accept write data
       -- Write Response channel (B)
   S_AXI_BREADY          : in std_logic;                                         -- Master ready to receive write response
   S_AXI_BRESP           : out std_logic_vector(1 downto 0);                     -- Write response from slave (OKAY or ERROR)
   S_AXI_BVALID          : out std_logic;                                        -- Slave asserts when write response is valid
       --Read Address channel (AR)
   S_AXI_ARADDR          : in std_logic_vector(G_ADDR_WIDTH-1 downto 0);         -- Read address from master to slave
   S_AXI_ARVALID         : in std_logic;                                         -- Master asserts when read address is valid
   S_AXI_ARREADY         : out std_logic;                                        -- Slave ready to accept read address
       -- Read channel (R)
   S_AXI_RREADY          : in std_logic;                                         -- Master ready to receive read data
   S_AXI_RDATA           : out std_logic_vector(G_DATA_WIDTH-1 downto 0);        -- Read data from slave to master
   S_AXI_RRESP           : out std_logic_vector(1 downto 0);                     -- Read response (OKAY or ERROR)
   S_AXI_RVALID          : out std_logic;                                        -- Slave asserts when read data is valid

   -- LANE + PHY interface
   ---------------------------------------
   -- to the LANE
   LANE_START            : out std_logic;                                        -- SpaceFibre lane start initialization signal
   AUTOSTART             : out std_logic;                                        -- Enables communication lane to initialize automatically when a link is established
   LANE_RESET            : out std_logic;                                        -- Reset Lane layer signal
   PARALLEL_LOOPBACK_EN  : out std_logic;                                        -- Parallel loopback enables signal
   STANDBY_REASON        : out std_logic_vector(C_STDBYREASON_WIDTH-1 downto 0); -- Standby reason field

   -- to the PHY
   NEAR_END_SERIAL_LB_EN : out std_logic;                                        -- Near-End Serial Loopback
   FAR_END_SERIAL_LB_EN  : out std_logic;                                        -- Far -End Serial Loopback

   -- from the LANE
   LANE_STATE            : in std_logic_vector(C_LANESTATE_WIDTH-1 downto 0);    -- Lane state field
   RX_ERROR_CNT          : in std_logic_vector(C_RX_ERR_CNT_WIDTH-1 downto 0);   -- RX Error Counter
   RX_ERROR_OVF          : in std_logic;                                         -- RX Error Overflow
   LOSS_SIGNAL           : in std_logic;                                         -- Far-end lost Signal
   FAR_END_CAPA          : in std_logic_vector(C_FAR_CAPA_WIDTH-1 downto 0);     -- Far-end Capablities
   RX_POLARITY           : in std_logic;                                         -- RX Polarity

   -- to the DUT
   RST_DUT_N             : out std_logic                                         -- Reset DUT (active low)
   );
end LANE_CONFIGURATOR;

------------------------------------------------------------------------------------------------------------------
--                                                  ARCHITECTURE                                                --
------------------------------------------------------------------------------------------------------------------
architecture rtl of LANE_CONFIGURATOR is
---------------------------------------
-- TYPES
---------------------------------------
   type axi_wr_state_t is (IDLE_WAIT_WR_ADDR, WR_RESPONSE);                      -- Write states for FSM declaration
   type axi_rd_state_t is (IDLE_WAIT_RD_ADDR, RD_RESPONSE);                      -- Read states for FSM declaration

---------------------------------------
-- SIGNAL DECLARATION
---------------------------------------
   signal axi_wr_state : axi_wr_state_t;
   signal axi_rd_state : axi_rd_state_t;
   -- Registers
   ------------
   signal reg_lane_param   : std_logic_vector(G_DATA_WIDTH-1 downto 0);          -- Lane parameters register
   signal reg_lane_status  : std_logic_vector(G_DATA_WIDTH-1 downto 0);          -- Lane status register
   signal reg_phy_param    : std_logic_vector(G_DATA_WIDTH-1 downto 0);          -- PHY parameters register
   signal reg_global       : std_logic_vector(G_DATA_WIDTH-1 downto 0);          -- Global register
   -- internal signals
   ------------
   signal lane_start_pulse : std_logic;                                          -- SpaceFibre lane start initialization signal pulsed

   signal lane_state_i     : std_logic_vector(C_LANESTATE_WIDTH-1 downto 0);    -- Lane state field
   signal rx_error_cnt_i   : std_logic_vector(C_RX_ERR_CNT_WIDTH-1 downto 0);   -- RX Error Counter
   signal rx_error_ovf_i   : std_logic;                                         -- RX Error Overflow
   signal loss_signal_i    : std_logic;                                         -- Far-end lost Signal
   signal far_end_capa_i   : std_logic_vector(C_FAR_CAPA_WIDTH-1 downto 0);     -- Far-end Capablities
   signal rx_polarity_i    : std_logic;                                         -- RX Polarity
   -- inputs resynchronization
   signal outputs_to_sync  : std_logic_vector(13 downto 0);
   signal outputs_to_dut   : std_logic_vector(13 downto 0);
   -- inputs resynchronization
   signal inputs_to_sync   : std_logic_vector(22 downto 0);
   signal inputs_to_model  : std_logic_vector(22 downto 0);
   begin
---------------------------------------
-- SIGNAL CONNECTION
---------------------------------------
   outputs_to_sync(0)           <= reg_lane_param(C_LANESTART_BTFD) or lane_start_pulse;
   outputs_to_sync(1)           <= reg_lane_param(C_AUTOSTART_BTFD);
   outputs_to_sync(2)           <= reg_lane_param(C_LANERESET_BTFD);
   outputs_to_sync(3)           <= reg_lane_param(C_PARALLEL_LPB_BTFD);
   outputs_to_sync(11 downto 4) <= reg_lane_param(C_STDBREASON_MAX_BTFD downto C_PARALLEL_LPB_BTFD +1);
   outputs_to_sync(12)          <= reg_phy_param(C_NEAR_END_LPB_BTFD);
   outputs_to_sync(13)          <= reg_phy_param(C_FAR_END_LPB_BTFD);

   LANE_START                   <= outputs_to_dut(0);
   AUTOSTART                    <= outputs_to_dut(1);
   LANE_RESET                   <= outputs_to_dut(2);
   PARALLEL_LOOPBACK_EN         <= outputs_to_dut(3);
   STANDBY_REASON               <= outputs_to_dut(11 downto 4);
   NEAR_END_SERIAL_LB_EN        <= outputs_to_dut(12);
   FAR_END_SERIAL_LB_EN         <= outputs_to_dut(13);

   inputs_to_sync(3 downto 0)   <= LANE_STATE;
   inputs_to_sync(11 downto 4)  <= RX_ERROR_CNT;
   inputs_to_sync(12)           <= RX_ERROR_OVF;
   inputs_to_sync(13)           <= LOSS_SIGNAL;
   inputs_to_sync(21 downto 14) <= FAR_END_CAPA;
   inputs_to_sync(22)           <= RX_POLARITY;

   lane_state_i                 <= inputs_to_model(3 downto 0);
   rx_error_cnt_i               <= inputs_to_model(11 downto 4);
   rx_error_ovf_i               <= inputs_to_model(12);
   loss_signal_i                <= inputs_to_model(13);
   far_end_capa_i               <= inputs_to_model(21 downto 14);
   rx_polarity_i                <= inputs_to_model(22);

   lane_start_pulse             <= reg_lane_param(C_LANESTART_PULSE_BTFD);
   RST_DUT_N                    <= reg_global(C_RST_DUT_BTFD);

---------------------------------------
-- INSTANCIATION
---------------------------------------
  ---------------------------------------------------------------------------
  -- INSTANCE: I_RESYNC_OUT
  -- Description : Resynchronize signals from the model at CLK to the CLK_TX clock
  ---------------------------------------------------------------------------
  I_RESYNC_OUT: entity work.resync_double
  generic map (
   VECTOR_SIZE => outputs_to_sync'length
  )
  port map (
   -- system signals
   clk    => CLK_TX,                                                               --- main clock
   rst_n  => RST_TXCLK_N,                                                          --- main reset (active low)
   -- I/Os
   input  => outputs_to_sync,                                                      --- vector to synchronize
   output => outputs_to_dut                                                        --- double synchronized vector
  );
  ---------------------------------------------------------------------------
  -- INSTANCE: I_RESYNC_IN
  -- Description : Resynchronize signals from the DUT at CLK_TX to the CLK clock
   ---------------------------------------------------------------------------
  I_RESYNC_IN: entity work.resync_double
  generic map (
   VECTOR_SIZE => inputs_to_sync'length
  )
  port map (
   -- system signals
   clk    => CLK,                                                                  --- main clock
   rst_n  => RST_N,                                                                --- main reset (active low)
   -- I/Os
   input  => inputs_to_sync,                                                       --- vector to synchronize
   output => inputs_to_model                                                       --- double synchronized vector
  );
---------------------------------------
-- PROCESS
---------------------------------------
   ---------------------------------------------------------------------------
   -- PROCESS: P_AXI_READ
   -- Description : AXI4 Lite reading process
   ---------------------------------------------------------------------------
   P_AXI_READ : process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N ='0') then
         axi_rd_state    <= IDLE_WAIT_RD_ADDR;
         S_AXI_ARREADY   <= '1';               -- Ready for new request
         S_AXI_RRESP     <= "00";              -- OKAY default response
         S_AXI_RDATA     <= (others => '0');   -- Default data at zero
         S_AXI_RVALID    <= '0';               -- Default read validity at zero
      elsif rising_edge(CLK) then
         case axi_rd_state is
            -- Waiting for a read request
            when IDLE_WAIT_RD_ADDR =>
               S_AXI_ARREADY <= '1';     -- Ready for new read request
               if (S_AXI_ARVALID = '1') then
                   S_AXI_ARREADY <= '0'; -- Ready signal deasserted to indicate request processing
                   -- Parameters lane register address
                   if (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_LANE_PARAM) then
                       S_AXI_RDATA  <= reg_lane_param;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Status lane register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_LANE_STATUS) then
                       S_AXI_RDATA  <= reg_lane_status;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Parameters PHY register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_PHY_PARAM) then
                       S_AXI_RDATA  <= reg_phy_param;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_GLOBAL) then
                       S_AXI_RDATA  <= reg_global;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Unrecognized address
                   else
                       S_AXI_RDATA  <= (others => '0');   -- Default response data
                       S_AXI_RRESP  <= "10";              -- Error response (SLVERR)
                       S_AXI_RVALID <= '1';               -- Response valid
                       axi_rd_state <= RD_RESPONSE;       -- Send the error response
                   end if;
               -- No read request received
               else
                   axi_rd_state <= IDLE_WAIT_RD_ADDR;
               end if;
            -- Responding to the read request
            when RD_RESPONSE =>
               -- Waiting for data reception confirmation from the master
               if (S_AXI_RREADY = '1') then
                   S_AXI_RVALID  <= '0';               -- Deassertion of response validity
                   S_AXI_RDATA   <= (others => '0');   -- Data reset
                   S_AXI_RRESP   <= "00";              -- Default OKAY response
                   axi_rd_state <= IDLE_WAIT_RD_ADDR;
               -- Wait until the master's reception confirmation is received
               else
                   axi_rd_state <= RD_RESPONSE;
               end if;
            -- Unrecognized state, return to IDLE state
            when others =>
               axi_rd_state <= IDLE_WAIT_RD_ADDR;
         end case;
      end if;
   end process P_AXI_READ;
   ---------------------------------------------------------------------------
   -- PROCESS: P_AXI_WRITE
   -- Description : AXI4 Lite writing process
   ---------------------------------------------------------------------------
   P_AXI_WRITE: process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N = '0') then
         axi_wr_state    <= IDLE_WAIT_WR_ADDR;
         S_AXI_AWREADY   <= '1';                 -- Ready for new request
         S_AXI_WREADY    <= '1';                 -- Ready to receive write data
         S_AXI_BRESP     <= "00";                -- OKAY default response
         S_AXI_BVALID    <= '0';                 -- Default write response validity
         reg_lane_param  <= init_lc_lane_param;
         reg_phy_param   <= init_lc_phy_param;
         reg_global      <= init_lc_global;
      elsif rising_edge(CLK) then
         if (lane_start_pulse ='1') then
            reg_lane_param(C_LANESTART_PULSE_BTFD)  <= '0';  -- Reset model start bit
         end if;
         case axi_wr_state is
            -- Waiting for a write request
            when IDLE_WAIT_WR_ADDR =>
               S_AXI_AWREADY   <= '1';              -- Ready for new request
               S_AXI_WREADY     <= '1';
               if (S_AXI_AWVALID = '1' and S_AXI_WVALID ='1') then
                  S_AXI_AWREADY   <= '0';           -- Ready signals deasserted to indicate request processing
                  S_AXI_WREADY    <= '0';
                  -- Parameters lane register address
                  if (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_LANE_PARAM) then
                     reg_lane_param <= S_AXI_WDATA; -- Write lane parameters
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Parameters phy register address
                  elsif (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_PHY_PARAM) then
                     reg_phy_param  <= S_AXI_WDATA; -- Write phy parameters
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  elsif (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_LC_GLOBAL) then
                     reg_global     <= S_AXI_WDATA; -- Write global signals
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Unrecognized address
                  else
                     S_AXI_BRESP  <= "10";          -- Error response (SLVERR)
                     S_AXI_BVALID <= '1';           -- Response valid
                     axi_wr_state <= WR_RESPONSE;
                  end if;
               -- No write request received
               else
                  axi_wr_state <= IDLE_WAIT_WR_ADDR;
               end if;
            -- Responding to the write request
            when WR_RESPONSE =>
               -- Waiting for response reception confirmation from the master
               if (S_AXI_BREADY  = '1') then
                  S_AXI_BVALID    <= '0';           -- Reset response validity
                  S_AXI_BRESP     <= "00";          -- Default OKAY response
                  axi_wr_state <= IDLE_WAIT_WR_ADDR;
               -- Wait until the master's reception confirmation is received
               else
                  axi_wr_state <= WR_RESPONSE;
               end if;
            -- Unrecognized state, return to IDLE state
            when others =>
                axi_wr_state <= IDLE_WAIT_WR_ADDR;
         end case;
      end if;
   end process P_AXI_WRITE;
   ---------------------------------------------------------------------------
   -- PROCESS: P_STATUS
   -- Description : update status register
   ---------------------------------------------------------------------------
   P_STATUS : process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N ='0') then
         reg_lane_status                                                      <= (others => '0');
      elsif rising_edge(CLK) then
         reg_lane_status(C_RX_POLARITY_BTFD)                                  <= rx_polarity_i;
         reg_lane_status(C_FAR_CAPA_MAX_BTFD downto C_FAR_LOST_SIG_BTFD+1)    <= far_end_capa_i;
         reg_lane_status(C_FAR_LOST_SIG_BTFD)                                 <= loss_signal_i;
         reg_lane_status(C_RX_ERR_OVF_BTFD)                                   <= rx_error_ovf_i;
         reg_lane_status(C_RX_ERR_CNT_MAX_BTFD downto C_LANESTATE_MAX_BTFD+1) <= rx_error_cnt_i;
         reg_lane_status(C_LANESTATE_MAX_BTFD downto 0)                       <= lane_state_i;
      end if;
   end process P_STATUS;
end rtl;
