`include "B_DSP_OUTPUT58_TEST_defines.vh"

reg [`DSP_OUTPUT58_TEST_DATA_SZ-1:0] ATTR [0:`DSP_OUTPUT58_TEST_ADDR_N-1];
reg [120:1] AUTORESET_PATDET_REG = AUTORESET_PATDET;
reg [40:1] AUTORESET_PRIORITY_REG = AUTORESET_PRIORITY;
reg [48:1] DSP_MODE_REG = DSP_MODE;
reg [56:1] EN_SCAN_REG = EN_SCAN;
reg IS_RSTP_INVERTED_REG = IS_RSTP_INVERTED;
reg [40:1] LEGACY_REG = LEGACY;
reg [31:0] PREG_REG = PREG;
reg [40:1] RESET_MODE_REG = RESET_MODE;

initial begin
  ATTR[`DSP_OUTPUT58_TEST__AUTORESET_PATDET] = AUTORESET_PATDET;
  ATTR[`DSP_OUTPUT58_TEST__AUTORESET_PRIORITY] = AUTORESET_PRIORITY;
  ATTR[`DSP_OUTPUT58_TEST__DSP_MODE] = DSP_MODE;
  ATTR[`DSP_OUTPUT58_TEST__EN_SCAN] = EN_SCAN;
  ATTR[`DSP_OUTPUT58_TEST__IS_RSTP_INVERTED] = IS_RSTP_INVERTED;
  ATTR[`DSP_OUTPUT58_TEST__LEGACY] = LEGACY;
  ATTR[`DSP_OUTPUT58_TEST__PREG] = PREG;
  ATTR[`DSP_OUTPUT58_TEST__RESET_MODE] = RESET_MODE;
end

always @(trig_attr) begin
  AUTORESET_PATDET_REG = ATTR[`DSP_OUTPUT58_TEST__AUTORESET_PATDET];
  AUTORESET_PRIORITY_REG = ATTR[`DSP_OUTPUT58_TEST__AUTORESET_PRIORITY];
  DSP_MODE_REG = ATTR[`DSP_OUTPUT58_TEST__DSP_MODE];
  EN_SCAN_REG = ATTR[`DSP_OUTPUT58_TEST__EN_SCAN];
  IS_RSTP_INVERTED_REG = ATTR[`DSP_OUTPUT58_TEST__IS_RSTP_INVERTED];
  LEGACY_REG = ATTR[`DSP_OUTPUT58_TEST__LEGACY];
  PREG_REG = ATTR[`DSP_OUTPUT58_TEST__PREG];
  RESET_MODE_REG = ATTR[`DSP_OUTPUT58_TEST__RESET_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_OUTPUT58_TEST_ADDR_SZ-1:0] addr;
  input  [`DSP_OUTPUT58_TEST_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_OUTPUT58_TEST_DATA_SZ-1:0] read_attr;
  input  [`DSP_OUTPUT58_TEST_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
