// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IBUFDS_DIFF_OUT_IBUFDISABLE_DEFINES_VH
`else
`define B_IBUFDS_DIFF_OUT_IBUFDISABLE_DEFINES_VH

// Look-up table parameters
//

`define IBUFDS_DIFF_OUT_IBUFDISABLE_ADDR_N  6
`define IBUFDS_DIFF_OUT_IBUFDISABLE_ADDR_SZ 32
`define IBUFDS_DIFF_OUT_IBUFDISABLE_DATA_SZ 144

// Attribute addresses
//

`define IBUFDS_DIFF_OUT_IBUFDISABLE__DIFF_TERM    32'h00000000
`define IBUFDS_DIFF_OUT_IBUFDISABLE__DIFF_TERM_SZ 40

`define IBUFDS_DIFF_OUT_IBUFDISABLE__DQS_BIAS    32'h00000001
`define IBUFDS_DIFF_OUT_IBUFDISABLE__DQS_BIAS_SZ 40

`define IBUFDS_DIFF_OUT_IBUFDISABLE__IBUF_LOW_PWR    32'h00000002
`define IBUFDS_DIFF_OUT_IBUFDISABLE__IBUF_LOW_PWR_SZ 40

`define IBUFDS_DIFF_OUT_IBUFDISABLE__IOSTANDARD    32'h00000003
`define IBUFDS_DIFF_OUT_IBUFDISABLE__IOSTANDARD_SZ 56

`define IBUFDS_DIFF_OUT_IBUFDISABLE__SIM_DEVICE    32'h00000004
`define IBUFDS_DIFF_OUT_IBUFDISABLE__SIM_DEVICE_SZ 144

`define IBUFDS_DIFF_OUT_IBUFDISABLE__USE_IBUFDISABLE    32'h00000005
`define IBUFDS_DIFF_OUT_IBUFDISABLE__USE_IBUFDISABLE_SZ 72

`endif  // B_IBUFDS_DIFF_OUT_IBUFDISABLE_DEFINES_VH