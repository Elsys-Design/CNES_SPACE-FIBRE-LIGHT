-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description :
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
  use phy_plus_lane_lib.all;
  use phy_plus_lane_lib.pkg_phy_plus_lane.all;

entity lane_ctrl_word_detect is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP

      -- RX control flag signals to from lane_init fsm
      NO_SIGNAL                        : out std_logic;                       --! Flag no signal are received
      RX_NEW_WORD                      : out std_logic;                       --! Flag new word has been received
      DETECTED_INIT1                   : out std_logic;                       --! Flag INIT1 control word rxed
      DETECTED_INIT2                   : out std_logic;                       --! Flag INIT2 control word rxed
      DETECTED_INIT3                   : out std_logic;                       --! Flag INIT3 control word rxed
      DETECTED_INV_INIT1               : out std_logic;                       --! Flag INV_INIT1 control word rxed
      DETECTED_INV_INIT2               : out std_logic;                       --! Flag INV_INIT2 control word rxed
      DETECTED_RXERR_WORD              : out std_logic;                       --! Flag RXERR detected
      DETECTED_LOSS_SIGNAL             : out std_logic;                       --! Flag LOSS_SIGNAL detected
      DETECTED_STANDBY                 : out std_logic;                       --! Flag STANDBY detected
      COMMA_K287_RXED                  : out std_logic;                       --! Flag Comma K28.7 has been received
      CAPABILITY                       : out std_logic_vector(07 downto 00);  --! Capability from INIT3 control word (31 downto 24)
      SEND_RXERR                       : in  std_logic;                       --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
      NO_SIGNAL_DETECTION_ENABLED      : in  std_logic;                       --! Flag to enable the no signal function
      ENABLE_TRANSM_DATA               : in  std_logic;                       --! Flag to enable the transmision of data

      -- RX signal from rx_sync_fsm/parallel_loopback
      DATA_RX_FROM_RSF                 : in  std_logic_vector(31 downto 00);  --! 32-bit data from rx_sync_fsm
      VALID_K_CARAC_FROM_RSF           : in  std_logic_vector(03 downto 00);  --! 4-bit valid K character flags from rx_sync_fsm
      DATA_RDY_FROM_RSF                : in  std_logic;                       --! Data valid flag from rx_sync_fsm

      -- RX signals to DATA-LINK
      DATA_RX_TO_DL                    : out std_logic_vector(31 downto 00);  --! 32-bit data to Data-link layer
      VALID_K_CARAC_TO_DL              : out std_logic_vector(03 downto 00);  --! 4-bit valid K character flags to Data-link layer
      DATA_RDY_TO_DL                   : out std_logic                        --! Data valid flag to Data-link layer
   );
end lane_ctrl_word_detect;

architecture rtl of lane_ctrl_word_detect is
----------------------------- Declaration signals -----------------------------
signal data_rx_to_dl_i                 : std_logic_vector(31 downto 00);      --! 32-bit data to Data-link layer
signal valid_k_charac_to_dl_i          : std_logic_vector(03 downto 00);      --! 4-bit valid K character flags to Data-link layer
signal data_rdy_to_dl_i                : std_logic;                           --! Data valid flag to Data-link layer
signal enable_transm_data_r            : std_logic;                           --! Transmission of data flag from init FSM
signal enable_transm_data_rr           : std_logic;                           --! Transmission of data flag from init FSM

begin

-- Detection of the control words
   p_ctrl_word_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         RX_NEW_WORD             <= '0';
         DETECTED_INIT1          <= '0';
         DETECTED_INIT2          <= '0';
         DETECTED_INIT3          <= '0';
         DETECTED_INV_INIT1      <= '0';
         DETECTED_INV_INIT2      <= '0';
         COMMA_K287_RXED         <= '0';
         DETECTED_LOSS_SIGNAL    <= '0';
         DETECTED_STANDBY        <= '0';
         data_rx_to_dl_i         <= (others => '0');
         valid_k_charac_to_dl_i  <= (others => '0');
         data_rdy_to_dl_i        <= '0';
         DETECTED_RXERR_WORD     <= '0';
         CAPABILITY              <= (others => '0');
         enable_transm_data_r    <= '0';

      elsif rising_edge(CLK) then
         
         enable_transm_data_r <= ENABLE_TRANSM_DATA;
         enable_transm_data_rr <= enable_transm_data_r;
         if DATA_RDY_FROM_RSF = '1' then                                   -- When new data is received

            if DATA_RX_FROM_RSF = C_INIT1_WORD and VALID_K_CARAC_FROM_RSF = "0001" then                        -- INIT1 control word detected
               DETECTED_INIT1          <= '1';                             -- Set INIT1 flag detected to '1'
               RX_NEW_WORD             <= '1';
            elsif DATA_RX_FROM_RSF = C_INIT2_WORD and VALID_K_CARAC_FROM_RSF = "0001" then                     -- INIT2 control word detected
               DETECTED_INIT2          <= '1';                             -- Set INIT2 flag detected to '1'
               RX_NEW_WORD             <= '1';
            elsif DATA_RX_FROM_RSF(23 downto 00) = C_INIT3_WORD and VALID_K_CARAC_FROM_RSF = "0001" then       -- INIT3 control word detected
               DETECTED_INIT3          <= '1';                             -- Set INIT3 flag detected to '1'
               RX_NEW_WORD             <= '1';
               CAPABILITY              <= DATA_RX_FROM_RSF(31 downto 24);
            elsif DATA_RX_FROM_RSF = C_I_INIT1_WORD and VALID_K_CARAC_FROM_RSF = "0001" then                   -- INIT1 inversed control word detected
               DETECTED_INV_INIT1      <= '1';                             -- Set INIT1 inversed flag detected to '1'
               RX_NEW_WORD             <= '1';
            elsif DATA_RX_FROM_RSF = C_I_INIT2_WORD and VALID_K_CARAC_FROM_RSF = "0001" then                   -- INIT2 inversed control word detected
               DETECTED_INV_INIT2      <= '1';                             -- Set INIT2 inversed flag detected to '1'
               RX_NEW_WORD             <= '1';
            elsif DATA_RX_FROM_RSF(23 downto 00) = C_LOST_SIG_WORD and VALID_K_CARAC_FROM_RSF = "0001" then    -- LOST_SIGNAL control word detected
               DETECTED_LOSS_SIGNAL    <= '1';                             -- Set LOSS_SIGNAL detected flag to '1'
               COMMA_K287_RXED         <= '1';                             -- Set Comma 28.7 detected flag to '1'
               RX_NEW_WORD             <= '1';
            elsif DATA_RX_FROM_RSF(23 downto 00) = C_STANDBY_WORD and VALID_K_CARAC_FROM_RSF = "0001" then     -- STANDBY control word detected
               DETECTED_STANDBY        <= '1';                             -- Set STANDBY detected flag to '1'
               COMMA_K287_RXED         <= '1';                             -- Set Comma 28.7 detected flag to '1'
               RX_NEW_WORD             <= '1';
            elsif SEND_RXERR = '1' and VALID_K_CARAC_FROM_RSF = "0001" then                                    -- When lane_init_fsm get out from ACTIVE_ST
               data_rx_to_dl_i         <= C_RXERR_WORD;                    -- Send a RXERR control word to DATA-LINK layer
               valid_k_charac_to_dl_i  <= x"1";
               data_rdy_to_dl_i        <= '1';
            elsif enable_transm_data_rr = '1' and not((DATA_RX_FROM_RSF = C_IDLE_WORD or DATA_RX_FROM_RSF = C_SKIP_WORD) and VALID_K_CARAC_FROM_RSF = "0001") then
               data_rx_to_dl_i         <= DATA_RX_FROM_RSF;                -- Else transmit data received from IP to DATA_LINK layer
               valid_k_charac_to_dl_i  <= VALID_K_CARAC_FROM_RSF;
               data_rdy_to_dl_i        <= DATA_RDY_FROM_RSF;
               RX_NEW_WORD             <= '1';
               
               if DATA_RX_FROM_RSF = C_RXERR_WORD and VALID_K_CARAC_FROM_RSF = "0001" then
                  DETECTED_RXERR_WORD  <= '1';
               else
                  DETECTED_RXERR_WORD  <= '0';
               end if;
               -- reset all flags
               DETECTED_INIT1          <= '0';
               DETECTED_INIT2          <= '0';
               DETECTED_INIT3          <= '0';
               DETECTED_INV_INIT1      <= '0';
               DETECTED_INV_INIT2      <= '0';
               COMMA_K287_RXED         <= '0';
               DETECTED_LOSS_SIGNAL    <= '0';
               DETECTED_STANDBY        <= '0';
            elsif (DATA_RX_FROM_RSF = C_IDLE_WORD or DATA_RX_FROM_RSF = C_SKIP_WORD) and VALID_K_CARAC_FROM_RSF = "0001" then                      -- IDLE or SKIP control word detected
               COMMA_K287_RXED         <= '1';                             -- Set Comma 28.7 detected flag to '1'
               RX_NEW_WORD             <= '1';
               data_rx_to_dl_i         <= (others => '0');                -- Else transmit data received from IP to DATA_LINK layer
               valid_k_charac_to_dl_i  <= (others => '0');
               data_rdy_to_dl_i        <= '0';
               if DATA_RX_FROM_RSF = C_RXERR_WORD and VALID_K_CARAC_FROM_RSF = "0001" then
                  DETECTED_RXERR_WORD  <= '1';
               else
                  DETECTED_RXERR_WORD  <= '0';
               end if;
                                              -- reset all flags
               DETECTED_INIT1          <= '0';
               DETECTED_INIT2          <= '0';
               DETECTED_INIT3          <= '0';
               DETECTED_INV_INIT1      <= '0';
               DETECTED_INV_INIT2      <= '0';
               DETECTED_LOSS_SIGNAL    <= '0';
               DETECTED_STANDBY        <= '0';
            else
               data_rx_to_dl_i         <= (others => '0');                -- Else transmit data received from IP to DATA_LINK layer
               valid_k_charac_to_dl_i  <= (others => '0');
               data_rdy_to_dl_i        <= '0';
               RX_NEW_WORD             <= '1'; 

               if DATA_RX_FROM_RSF = C_RXERR_WORD and VALID_K_CARAC_FROM_RSF = "0001" then
                  DETECTED_RXERR_WORD  <= '1';
               else
                  DETECTED_RXERR_WORD  <= '0';
               end if;
                                              -- reset all flags
               DETECTED_INIT1          <= '0';
               DETECTED_INIT2          <= '0';
               DETECTED_INIT3          <= '0';
               DETECTED_INV_INIT1      <= '0';
               DETECTED_INV_INIT2      <= '0';
               COMMA_K287_RXED         <= '0';
               DETECTED_LOSS_SIGNAL    <= '0';
               DETECTED_STANDBY        <= '0';
            end if;

         else
            RX_NEW_WORD             <= '0';                                -- else reset all flags
            DETECTED_INIT1          <= '0';
            DETECTED_INIT2          <= '0';
            DETECTED_INIT3          <= '0';
            DETECTED_INV_INIT1      <= '0';
            DETECTED_INV_INIT2      <= '0';
            COMMA_K287_RXED         <= '0';
            DETECTED_LOSS_SIGNAL    <= '0';
            DETECTED_STANDBY        <= '0';
            data_rx_to_dl_i         <= (others => '0');
            valid_k_charac_to_dl_i  <= (others => '0');
            data_rdy_to_dl_i        <= '0';
            DETECTED_RXERR_WORD     <= '0';
         end if;

      end if;
   end process p_ctrl_word_detection;




   p_no_signal_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         NO_SIGNAL   <= '0';
      elsif rising_edge(CLK) then

         if NO_SIGNAL_DETECTION_ENABLED = '1' then
            NO_SIGNAL   <= '0';
         else
            NO_SIGNAL   <= '0';
         end if;
      end if;
   end process p_no_signal_detection;

-- Outputs
DATA_RX_TO_DL         <= data_rx_to_dl_i;
VALID_K_CARAC_TO_DL   <= valid_k_charac_to_dl_i;
DATA_RDY_TO_DL        <= data_rdy_to_dl_i;

end architecture rtl;
