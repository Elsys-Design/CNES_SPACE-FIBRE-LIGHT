// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTF_CHANNEL_DEFINES_VH
`else
`define B_GTF_CHANNEL_DEFINES_VH

// Look-up table parameters
//

`define GTF_CHANNEL_ADDR_N  379
`define GTF_CHANNEL_ADDR_SZ 32
`define GTF_CHANNEL_DATA_SZ 88

// Attribute addresses
//

`define GTF_CHANNEL__ACJTAG_DEBUG_MODE    32'h00000000
`define GTF_CHANNEL__ACJTAG_DEBUG_MODE_SZ 1

`define GTF_CHANNEL__ACJTAG_MODE    32'h00000001
`define GTF_CHANNEL__ACJTAG_MODE_SZ 1

`define GTF_CHANNEL__ACJTAG_RESET    32'h00000002
`define GTF_CHANNEL__ACJTAG_RESET_SZ 1

`define GTF_CHANNEL__ADAPT_CFG0    32'h00000003
`define GTF_CHANNEL__ADAPT_CFG0_SZ 16

`define GTF_CHANNEL__ADAPT_CFG1    32'h00000004
`define GTF_CHANNEL__ADAPT_CFG1_SZ 16

`define GTF_CHANNEL__ADAPT_CFG2    32'h00000005
`define GTF_CHANNEL__ADAPT_CFG2_SZ 16

`define GTF_CHANNEL__A_RXOSCALRESET    32'h00000006
`define GTF_CHANNEL__A_RXOSCALRESET_SZ 1

`define GTF_CHANNEL__A_RXPROGDIVRESET    32'h00000007
`define GTF_CHANNEL__A_RXPROGDIVRESET_SZ 1

`define GTF_CHANNEL__A_RXTERMINATION    32'h00000008
`define GTF_CHANNEL__A_RXTERMINATION_SZ 1

`define GTF_CHANNEL__A_TXDIFFCTRL    32'h00000009
`define GTF_CHANNEL__A_TXDIFFCTRL_SZ 5

`define GTF_CHANNEL__A_TXPROGDIVRESET    32'h0000000a
`define GTF_CHANNEL__A_TXPROGDIVRESET_SZ 1

`define GTF_CHANNEL__CBCC_DATA_SOURCE_SEL    32'h0000000b
`define GTF_CHANNEL__CBCC_DATA_SOURCE_SEL_SZ 56

`define GTF_CHANNEL__CDR_SWAP_MODE_EN    32'h0000000c
`define GTF_CHANNEL__CDR_SWAP_MODE_EN_SZ 1

`define GTF_CHANNEL__CFOK_PWRSVE_EN    32'h0000000d
`define GTF_CHANNEL__CFOK_PWRSVE_EN_SZ 1

`define GTF_CHANNEL__CH_HSPMUX    32'h0000000e
`define GTF_CHANNEL__CH_HSPMUX_SZ 16

`define GTF_CHANNEL__CKCAL1_CFG_0    32'h0000000f
`define GTF_CHANNEL__CKCAL1_CFG_0_SZ 16

`define GTF_CHANNEL__CKCAL1_CFG_1    32'h00000010
`define GTF_CHANNEL__CKCAL1_CFG_1_SZ 16

`define GTF_CHANNEL__CKCAL1_CFG_2    32'h00000011
`define GTF_CHANNEL__CKCAL1_CFG_2_SZ 16

`define GTF_CHANNEL__CKCAL1_CFG_3    32'h00000012
`define GTF_CHANNEL__CKCAL1_CFG_3_SZ 16

`define GTF_CHANNEL__CKCAL2_CFG_0    32'h00000013
`define GTF_CHANNEL__CKCAL2_CFG_0_SZ 16

`define GTF_CHANNEL__CKCAL2_CFG_1    32'h00000014
`define GTF_CHANNEL__CKCAL2_CFG_1_SZ 16

`define GTF_CHANNEL__CKCAL2_CFG_2    32'h00000015
`define GTF_CHANNEL__CKCAL2_CFG_2_SZ 16

`define GTF_CHANNEL__CKCAL2_CFG_3    32'h00000016
`define GTF_CHANNEL__CKCAL2_CFG_3_SZ 16

`define GTF_CHANNEL__CKCAL2_CFG_4    32'h00000017
`define GTF_CHANNEL__CKCAL2_CFG_4_SZ 16

`define GTF_CHANNEL__CPLL_CFG0    32'h00000018
`define GTF_CHANNEL__CPLL_CFG0_SZ 16

`define GTF_CHANNEL__CPLL_CFG1    32'h00000019
`define GTF_CHANNEL__CPLL_CFG1_SZ 16

`define GTF_CHANNEL__CPLL_CFG2    32'h0000001a
`define GTF_CHANNEL__CPLL_CFG2_SZ 16

`define GTF_CHANNEL__CPLL_CFG3    32'h0000001b
`define GTF_CHANNEL__CPLL_CFG3_SZ 16

`define GTF_CHANNEL__CPLL_FBDIV    32'h0000001c
`define GTF_CHANNEL__CPLL_FBDIV_SZ 5

`define GTF_CHANNEL__CPLL_FBDIV_45    32'h0000001d
`define GTF_CHANNEL__CPLL_FBDIV_45_SZ 3

`define GTF_CHANNEL__CPLL_INIT_CFG0    32'h0000001e
`define GTF_CHANNEL__CPLL_INIT_CFG0_SZ 16

`define GTF_CHANNEL__CPLL_LOCK_CFG    32'h0000001f
`define GTF_CHANNEL__CPLL_LOCK_CFG_SZ 16

`define GTF_CHANNEL__CPLL_REFCLK_DIV    32'h00000020
`define GTF_CHANNEL__CPLL_REFCLK_DIV_SZ 5

`define GTF_CHANNEL__CTLE3_OCAP_EXT_CTRL    32'h00000021
`define GTF_CHANNEL__CTLE3_OCAP_EXT_CTRL_SZ 3

`define GTF_CHANNEL__CTLE3_OCAP_EXT_EN    32'h00000022
`define GTF_CHANNEL__CTLE3_OCAP_EXT_EN_SZ 1

`define GTF_CHANNEL__DDI_CTRL    32'h00000023
`define GTF_CHANNEL__DDI_CTRL_SZ 2

`define GTF_CHANNEL__DDI_REALIGN_WAIT    32'h00000024
`define GTF_CHANNEL__DDI_REALIGN_WAIT_SZ 5

`define GTF_CHANNEL__DELAY_ELEC    32'h00000025
`define GTF_CHANNEL__DELAY_ELEC_SZ 1

`define GTF_CHANNEL__DMONITOR_CFG0    32'h00000026
`define GTF_CHANNEL__DMONITOR_CFG0_SZ 10

`define GTF_CHANNEL__DMONITOR_CFG1    32'h00000027
`define GTF_CHANNEL__DMONITOR_CFG1_SZ 8

`define GTF_CHANNEL__ES_CLK_PHASE_SEL    32'h00000028
`define GTF_CHANNEL__ES_CLK_PHASE_SEL_SZ 1

`define GTF_CHANNEL__ES_CONTROL    32'h00000029
`define GTF_CHANNEL__ES_CONTROL_SZ 6

`define GTF_CHANNEL__ES_ERRDET_EN    32'h0000002a
`define GTF_CHANNEL__ES_ERRDET_EN_SZ 40

`define GTF_CHANNEL__ES_EYE_SCAN_EN    32'h0000002b
`define GTF_CHANNEL__ES_EYE_SCAN_EN_SZ 40

`define GTF_CHANNEL__ES_HORZ_OFFSET    32'h0000002c
`define GTF_CHANNEL__ES_HORZ_OFFSET_SZ 12

`define GTF_CHANNEL__ES_PRESCALE    32'h0000002d
`define GTF_CHANNEL__ES_PRESCALE_SZ 5

`define GTF_CHANNEL__ES_QUALIFIER0    32'h0000002e
`define GTF_CHANNEL__ES_QUALIFIER0_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER1    32'h0000002f
`define GTF_CHANNEL__ES_QUALIFIER1_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER2    32'h00000030
`define GTF_CHANNEL__ES_QUALIFIER2_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER3    32'h00000031
`define GTF_CHANNEL__ES_QUALIFIER3_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER4    32'h00000032
`define GTF_CHANNEL__ES_QUALIFIER4_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER5    32'h00000033
`define GTF_CHANNEL__ES_QUALIFIER5_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER6    32'h00000034
`define GTF_CHANNEL__ES_QUALIFIER6_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER7    32'h00000035
`define GTF_CHANNEL__ES_QUALIFIER7_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER8    32'h00000036
`define GTF_CHANNEL__ES_QUALIFIER8_SZ 16

`define GTF_CHANNEL__ES_QUALIFIER9    32'h00000037
`define GTF_CHANNEL__ES_QUALIFIER9_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK0    32'h00000038
`define GTF_CHANNEL__ES_QUAL_MASK0_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK1    32'h00000039
`define GTF_CHANNEL__ES_QUAL_MASK1_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK2    32'h0000003a
`define GTF_CHANNEL__ES_QUAL_MASK2_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK3    32'h0000003b
`define GTF_CHANNEL__ES_QUAL_MASK3_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK4    32'h0000003c
`define GTF_CHANNEL__ES_QUAL_MASK4_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK5    32'h0000003d
`define GTF_CHANNEL__ES_QUAL_MASK5_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK6    32'h0000003e
`define GTF_CHANNEL__ES_QUAL_MASK6_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK7    32'h0000003f
`define GTF_CHANNEL__ES_QUAL_MASK7_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK8    32'h00000040
`define GTF_CHANNEL__ES_QUAL_MASK8_SZ 16

`define GTF_CHANNEL__ES_QUAL_MASK9    32'h00000041
`define GTF_CHANNEL__ES_QUAL_MASK9_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK0    32'h00000042
`define GTF_CHANNEL__ES_SDATA_MASK0_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK1    32'h00000043
`define GTF_CHANNEL__ES_SDATA_MASK1_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK2    32'h00000044
`define GTF_CHANNEL__ES_SDATA_MASK2_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK3    32'h00000045
`define GTF_CHANNEL__ES_SDATA_MASK3_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK4    32'h00000046
`define GTF_CHANNEL__ES_SDATA_MASK4_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK5    32'h00000047
`define GTF_CHANNEL__ES_SDATA_MASK5_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK6    32'h00000048
`define GTF_CHANNEL__ES_SDATA_MASK6_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK7    32'h00000049
`define GTF_CHANNEL__ES_SDATA_MASK7_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK8    32'h0000004a
`define GTF_CHANNEL__ES_SDATA_MASK8_SZ 16

`define GTF_CHANNEL__ES_SDATA_MASK9    32'h0000004b
`define GTF_CHANNEL__ES_SDATA_MASK9_SZ 16

`define GTF_CHANNEL__EYESCAN_VP_RANGE    32'h0000004c
`define GTF_CHANNEL__EYESCAN_VP_RANGE_SZ 2

`define GTF_CHANNEL__EYE_SCAN_SWAP_EN    32'h0000004d
`define GTF_CHANNEL__EYE_SCAN_SWAP_EN_SZ 1

`define GTF_CHANNEL__FTS_DESKEW_SEQ_ENABLE    32'h0000004e
`define GTF_CHANNEL__FTS_DESKEW_SEQ_ENABLE_SZ 4

`define GTF_CHANNEL__FTS_LANE_DESKEW_CFG    32'h0000004f
`define GTF_CHANNEL__FTS_LANE_DESKEW_CFG_SZ 4

`define GTF_CHANNEL__FTS_LANE_DESKEW_EN    32'h00000050
`define GTF_CHANNEL__FTS_LANE_DESKEW_EN_SZ 40

`define GTF_CHANNEL__GEARBOX_MODE    32'h00000051
`define GTF_CHANNEL__GEARBOX_MODE_SZ 5

`define GTF_CHANNEL__ISCAN_CK_PH_SEL2    32'h00000052
`define GTF_CHANNEL__ISCAN_CK_PH_SEL2_SZ 1

`define GTF_CHANNEL__LOCAL_MASTER    32'h00000053
`define GTF_CHANNEL__LOCAL_MASTER_SZ 1

`define GTF_CHANNEL__LPBK_BIAS_CTRL    32'h00000054
`define GTF_CHANNEL__LPBK_BIAS_CTRL_SZ 3

`define GTF_CHANNEL__LPBK_EN_RCAL_B    32'h00000055
`define GTF_CHANNEL__LPBK_EN_RCAL_B_SZ 1

`define GTF_CHANNEL__LPBK_EXT_RCAL    32'h00000056
`define GTF_CHANNEL__LPBK_EXT_RCAL_SZ 4

`define GTF_CHANNEL__LPBK_IND_CTRL0    32'h00000057
`define GTF_CHANNEL__LPBK_IND_CTRL0_SZ 3

`define GTF_CHANNEL__LPBK_IND_CTRL1    32'h00000058
`define GTF_CHANNEL__LPBK_IND_CTRL1_SZ 3

`define GTF_CHANNEL__LPBK_IND_CTRL2    32'h00000059
`define GTF_CHANNEL__LPBK_IND_CTRL2_SZ 3

`define GTF_CHANNEL__LPBK_RG_CTRL    32'h0000005a
`define GTF_CHANNEL__LPBK_RG_CTRL_SZ 2

`define GTF_CHANNEL__MAC_CFG0    32'h0000005b
`define GTF_CHANNEL__MAC_CFG0_SZ 16

`define GTF_CHANNEL__MAC_CFG1    32'h0000005c
`define GTF_CHANNEL__MAC_CFG1_SZ 16

`define GTF_CHANNEL__MAC_CFG10    32'h0000005d
`define GTF_CHANNEL__MAC_CFG10_SZ 16

`define GTF_CHANNEL__MAC_CFG11    32'h0000005e
`define GTF_CHANNEL__MAC_CFG11_SZ 16

`define GTF_CHANNEL__MAC_CFG12    32'h0000005f
`define GTF_CHANNEL__MAC_CFG12_SZ 16

`define GTF_CHANNEL__MAC_CFG13    32'h00000060
`define GTF_CHANNEL__MAC_CFG13_SZ 16

`define GTF_CHANNEL__MAC_CFG14    32'h00000061
`define GTF_CHANNEL__MAC_CFG14_SZ 16

`define GTF_CHANNEL__MAC_CFG15    32'h00000062
`define GTF_CHANNEL__MAC_CFG15_SZ 16

`define GTF_CHANNEL__MAC_CFG2    32'h00000063
`define GTF_CHANNEL__MAC_CFG2_SZ 16

`define GTF_CHANNEL__MAC_CFG3    32'h00000064
`define GTF_CHANNEL__MAC_CFG3_SZ 16

`define GTF_CHANNEL__MAC_CFG4    32'h00000065
`define GTF_CHANNEL__MAC_CFG4_SZ 16

`define GTF_CHANNEL__MAC_CFG5    32'h00000066
`define GTF_CHANNEL__MAC_CFG5_SZ 16

`define GTF_CHANNEL__MAC_CFG6    32'h00000067
`define GTF_CHANNEL__MAC_CFG6_SZ 16

`define GTF_CHANNEL__MAC_CFG7    32'h00000068
`define GTF_CHANNEL__MAC_CFG7_SZ 16

`define GTF_CHANNEL__MAC_CFG8    32'h00000069
`define GTF_CHANNEL__MAC_CFG8_SZ 16

`define GTF_CHANNEL__MAC_CFG9    32'h0000006a
`define GTF_CHANNEL__MAC_CFG9_SZ 16

`define GTF_CHANNEL__PCS_RSVD0    32'h0000006b
`define GTF_CHANNEL__PCS_RSVD0_SZ 16

`define GTF_CHANNEL__PD_TRANS_TIME_FROM_P2    32'h0000006c
`define GTF_CHANNEL__PD_TRANS_TIME_FROM_P2_SZ 12

`define GTF_CHANNEL__PD_TRANS_TIME_NONE_P2    32'h0000006d
`define GTF_CHANNEL__PD_TRANS_TIME_NONE_P2_SZ 8

`define GTF_CHANNEL__PD_TRANS_TIME_TO_P2    32'h0000006e
`define GTF_CHANNEL__PD_TRANS_TIME_TO_P2_SZ 8

`define GTF_CHANNEL__PREIQ_FREQ_BST    32'h0000006f
`define GTF_CHANNEL__PREIQ_FREQ_BST_SZ 2

`define GTF_CHANNEL__RAW_MAC_CFG    32'h00000070
`define GTF_CHANNEL__RAW_MAC_CFG_SZ 16

`define GTF_CHANNEL__RCLK_SIPO_DLY_ENB    32'h00000071
`define GTF_CHANNEL__RCLK_SIPO_DLY_ENB_SZ 1

`define GTF_CHANNEL__RCLK_SIPO_INV_EN    32'h00000072
`define GTF_CHANNEL__RCLK_SIPO_INV_EN_SZ 1

`define GTF_CHANNEL__RCO_NEW_MAC_CFG0    32'h00000073
`define GTF_CHANNEL__RCO_NEW_MAC_CFG0_SZ 16

`define GTF_CHANNEL__RCO_NEW_MAC_CFG1    32'h00000074
`define GTF_CHANNEL__RCO_NEW_MAC_CFG1_SZ 16

`define GTF_CHANNEL__RCO_NEW_MAC_CFG2    32'h00000075
`define GTF_CHANNEL__RCO_NEW_MAC_CFG2_SZ 16

`define GTF_CHANNEL__RCO_NEW_MAC_CFG3    32'h00000076
`define GTF_CHANNEL__RCO_NEW_MAC_CFG3_SZ 16

`define GTF_CHANNEL__RCO_NEW_RAW_CFG0    32'h00000077
`define GTF_CHANNEL__RCO_NEW_RAW_CFG0_SZ 16

`define GTF_CHANNEL__RCO_NEW_RAW_CFG1    32'h00000078
`define GTF_CHANNEL__RCO_NEW_RAW_CFG1_SZ 16

`define GTF_CHANNEL__RCO_NEW_RAW_CFG2    32'h00000079
`define GTF_CHANNEL__RCO_NEW_RAW_CFG2_SZ 16

`define GTF_CHANNEL__RCO_NEW_RAW_CFG3    32'h0000007a
`define GTF_CHANNEL__RCO_NEW_RAW_CFG3_SZ 16

`define GTF_CHANNEL__RTX_BUF_CML_CTRL    32'h0000007b
`define GTF_CHANNEL__RTX_BUF_CML_CTRL_SZ 3

`define GTF_CHANNEL__RTX_BUF_TERM_CTRL    32'h0000007c
`define GTF_CHANNEL__RTX_BUF_TERM_CTRL_SZ 2

`define GTF_CHANNEL__RXBUFRESET_TIME    32'h0000007d
`define GTF_CHANNEL__RXBUFRESET_TIME_SZ 5

`define GTF_CHANNEL__RXBUF_EN    32'h0000007e
`define GTF_CHANNEL__RXBUF_EN_SZ 40

`define GTF_CHANNEL__RXCDRFREQRESET_TIME    32'h0000007f
`define GTF_CHANNEL__RXCDRFREQRESET_TIME_SZ 5

`define GTF_CHANNEL__RXCDRPHRESET_TIME    32'h00000080
`define GTF_CHANNEL__RXCDRPHRESET_TIME_SZ 5

`define GTF_CHANNEL__RXCDR_CFG0    32'h00000081
`define GTF_CHANNEL__RXCDR_CFG0_SZ 16

`define GTF_CHANNEL__RXCDR_CFG1    32'h00000082
`define GTF_CHANNEL__RXCDR_CFG1_SZ 16

`define GTF_CHANNEL__RXCDR_CFG2    32'h00000083
`define GTF_CHANNEL__RXCDR_CFG2_SZ 16

`define GTF_CHANNEL__RXCDR_CFG3    32'h00000084
`define GTF_CHANNEL__RXCDR_CFG3_SZ 16

`define GTF_CHANNEL__RXCDR_CFG4    32'h00000085
`define GTF_CHANNEL__RXCDR_CFG4_SZ 16

`define GTF_CHANNEL__RXCDR_CFG5    32'h00000086
`define GTF_CHANNEL__RXCDR_CFG5_SZ 16

`define GTF_CHANNEL__RXCDR_FR_RESET_ON_EIDLE    32'h00000087
`define GTF_CHANNEL__RXCDR_FR_RESET_ON_EIDLE_SZ 1

`define GTF_CHANNEL__RXCDR_HOLD_DURING_EIDLE    32'h00000088
`define GTF_CHANNEL__RXCDR_HOLD_DURING_EIDLE_SZ 1

`define GTF_CHANNEL__RXCDR_LOCK_CFG0    32'h00000089
`define GTF_CHANNEL__RXCDR_LOCK_CFG0_SZ 16

`define GTF_CHANNEL__RXCDR_LOCK_CFG1    32'h0000008a
`define GTF_CHANNEL__RXCDR_LOCK_CFG1_SZ 16

`define GTF_CHANNEL__RXCDR_LOCK_CFG2    32'h0000008b
`define GTF_CHANNEL__RXCDR_LOCK_CFG2_SZ 16

`define GTF_CHANNEL__RXCDR_LOCK_CFG3    32'h0000008c
`define GTF_CHANNEL__RXCDR_LOCK_CFG3_SZ 16

`define GTF_CHANNEL__RXCDR_LOCK_CFG4    32'h0000008d
`define GTF_CHANNEL__RXCDR_LOCK_CFG4_SZ 16

`define GTF_CHANNEL__RXCDR_PH_RESET_ON_EIDLE    32'h0000008e
`define GTF_CHANNEL__RXCDR_PH_RESET_ON_EIDLE_SZ 1

`define GTF_CHANNEL__RXCFOK_CFG0    32'h0000008f
`define GTF_CHANNEL__RXCFOK_CFG0_SZ 16

`define GTF_CHANNEL__RXCFOK_CFG1    32'h00000090
`define GTF_CHANNEL__RXCFOK_CFG1_SZ 16

`define GTF_CHANNEL__RXCFOK_CFG2    32'h00000091
`define GTF_CHANNEL__RXCFOK_CFG2_SZ 16

`define GTF_CHANNEL__RXCKCAL1_IQ_LOOP_RST_CFG    32'h00000092
`define GTF_CHANNEL__RXCKCAL1_IQ_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL1_I_LOOP_RST_CFG    32'h00000093
`define GTF_CHANNEL__RXCKCAL1_I_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL1_Q_LOOP_RST_CFG    32'h00000094
`define GTF_CHANNEL__RXCKCAL1_Q_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL2_DX_LOOP_RST_CFG    32'h00000095
`define GTF_CHANNEL__RXCKCAL2_DX_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL2_D_LOOP_RST_CFG    32'h00000096
`define GTF_CHANNEL__RXCKCAL2_D_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL2_S_LOOP_RST_CFG    32'h00000097
`define GTF_CHANNEL__RXCKCAL2_S_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXCKCAL2_X_LOOP_RST_CFG    32'h00000098
`define GTF_CHANNEL__RXCKCAL2_X_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__RXDFELPMRESET_TIME    32'h00000099
`define GTF_CHANNEL__RXDFELPMRESET_TIME_SZ 7

`define GTF_CHANNEL__RXDFELPM_KL_CFG0    32'h0000009a
`define GTF_CHANNEL__RXDFELPM_KL_CFG0_SZ 16

`define GTF_CHANNEL__RXDFELPM_KL_CFG1    32'h0000009b
`define GTF_CHANNEL__RXDFELPM_KL_CFG1_SZ 16

`define GTF_CHANNEL__RXDFELPM_KL_CFG2    32'h0000009c
`define GTF_CHANNEL__RXDFELPM_KL_CFG2_SZ 16

`define GTF_CHANNEL__RXDFE_CFG0    32'h0000009d
`define GTF_CHANNEL__RXDFE_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_CFG1    32'h0000009e
`define GTF_CHANNEL__RXDFE_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_GC_CFG0    32'h0000009f
`define GTF_CHANNEL__RXDFE_GC_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_GC_CFG1    32'h000000a0
`define GTF_CHANNEL__RXDFE_GC_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_GC_CFG2    32'h000000a1
`define GTF_CHANNEL__RXDFE_GC_CFG2_SZ 16

`define GTF_CHANNEL__RXDFE_H2_CFG0    32'h000000a2
`define GTF_CHANNEL__RXDFE_H2_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H2_CFG1    32'h000000a3
`define GTF_CHANNEL__RXDFE_H2_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H3_CFG0    32'h000000a4
`define GTF_CHANNEL__RXDFE_H3_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H3_CFG1    32'h000000a5
`define GTF_CHANNEL__RXDFE_H3_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H4_CFG0    32'h000000a6
`define GTF_CHANNEL__RXDFE_H4_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H4_CFG1    32'h000000a7
`define GTF_CHANNEL__RXDFE_H4_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H5_CFG0    32'h000000a8
`define GTF_CHANNEL__RXDFE_H5_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H5_CFG1    32'h000000a9
`define GTF_CHANNEL__RXDFE_H5_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H6_CFG0    32'h000000aa
`define GTF_CHANNEL__RXDFE_H6_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H6_CFG1    32'h000000ab
`define GTF_CHANNEL__RXDFE_H6_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H7_CFG0    32'h000000ac
`define GTF_CHANNEL__RXDFE_H7_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H7_CFG1    32'h000000ad
`define GTF_CHANNEL__RXDFE_H7_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H8_CFG0    32'h000000ae
`define GTF_CHANNEL__RXDFE_H8_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H8_CFG1    32'h000000af
`define GTF_CHANNEL__RXDFE_H8_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_H9_CFG0    32'h000000b0
`define GTF_CHANNEL__RXDFE_H9_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_H9_CFG1    32'h000000b1
`define GTF_CHANNEL__RXDFE_H9_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HA_CFG0    32'h000000b2
`define GTF_CHANNEL__RXDFE_HA_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HA_CFG1    32'h000000b3
`define GTF_CHANNEL__RXDFE_HA_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HB_CFG0    32'h000000b4
`define GTF_CHANNEL__RXDFE_HB_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HB_CFG1    32'h000000b5
`define GTF_CHANNEL__RXDFE_HB_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HC_CFG0    32'h000000b6
`define GTF_CHANNEL__RXDFE_HC_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HC_CFG1    32'h000000b7
`define GTF_CHANNEL__RXDFE_HC_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HD_CFG0    32'h000000b8
`define GTF_CHANNEL__RXDFE_HD_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HD_CFG1    32'h000000b9
`define GTF_CHANNEL__RXDFE_HD_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HE_CFG0    32'h000000ba
`define GTF_CHANNEL__RXDFE_HE_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HE_CFG1    32'h000000bb
`define GTF_CHANNEL__RXDFE_HE_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_HF_CFG0    32'h000000bc
`define GTF_CHANNEL__RXDFE_HF_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_HF_CFG1    32'h000000bd
`define GTF_CHANNEL__RXDFE_HF_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_KH_CFG0    32'h000000be
`define GTF_CHANNEL__RXDFE_KH_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_KH_CFG1    32'h000000bf
`define GTF_CHANNEL__RXDFE_KH_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_KH_CFG2    32'h000000c0
`define GTF_CHANNEL__RXDFE_KH_CFG2_SZ 16

`define GTF_CHANNEL__RXDFE_KH_CFG3    32'h000000c1
`define GTF_CHANNEL__RXDFE_KH_CFG3_SZ 16

`define GTF_CHANNEL__RXDFE_OS_CFG0    32'h000000c2
`define GTF_CHANNEL__RXDFE_OS_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_OS_CFG1    32'h000000c3
`define GTF_CHANNEL__RXDFE_OS_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_UT_CFG0    32'h000000c4
`define GTF_CHANNEL__RXDFE_UT_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_UT_CFG1    32'h000000c5
`define GTF_CHANNEL__RXDFE_UT_CFG1_SZ 16

`define GTF_CHANNEL__RXDFE_UT_CFG2    32'h000000c6
`define GTF_CHANNEL__RXDFE_UT_CFG2_SZ 16

`define GTF_CHANNEL__RXDFE_VP_CFG0    32'h000000c7
`define GTF_CHANNEL__RXDFE_VP_CFG0_SZ 16

`define GTF_CHANNEL__RXDFE_VP_CFG1    32'h000000c8
`define GTF_CHANNEL__RXDFE_VP_CFG1_SZ 16

`define GTF_CHANNEL__RXDLY_CFG    32'h000000c9
`define GTF_CHANNEL__RXDLY_CFG_SZ 16

`define GTF_CHANNEL__RXDLY_LCFG    32'h000000ca
`define GTF_CHANNEL__RXDLY_LCFG_SZ 16

`define GTF_CHANNEL__RXDLY_RAW_CFG    32'h000000cb
`define GTF_CHANNEL__RXDLY_RAW_CFG_SZ 16

`define GTF_CHANNEL__RXDLY_RAW_LCFG    32'h000000cc
`define GTF_CHANNEL__RXDLY_RAW_LCFG_SZ 16

`define GTF_CHANNEL__RXELECIDLE_CFG    32'h000000cd
`define GTF_CHANNEL__RXELECIDLE_CFG_SZ 72

`define GTF_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR    32'h000000ce
`define GTF_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR_SZ 3

`define GTF_CHANNEL__RXGEARBOX_EN    32'h000000cf
`define GTF_CHANNEL__RXGEARBOX_EN_SZ 40

`define GTF_CHANNEL__RXISCANRESET_TIME    32'h000000d0
`define GTF_CHANNEL__RXISCANRESET_TIME_SZ 5

`define GTF_CHANNEL__RXLPM_CFG    32'h000000d1
`define GTF_CHANNEL__RXLPM_CFG_SZ 16

`define GTF_CHANNEL__RXLPM_GC_CFG    32'h000000d2
`define GTF_CHANNEL__RXLPM_GC_CFG_SZ 16

`define GTF_CHANNEL__RXLPM_KH_CFG0    32'h000000d3
`define GTF_CHANNEL__RXLPM_KH_CFG0_SZ 16

`define GTF_CHANNEL__RXLPM_KH_CFG1    32'h000000d4
`define GTF_CHANNEL__RXLPM_KH_CFG1_SZ 16

`define GTF_CHANNEL__RXLPM_OS_CFG0    32'h000000d5
`define GTF_CHANNEL__RXLPM_OS_CFG0_SZ 16

`define GTF_CHANNEL__RXLPM_OS_CFG1    32'h000000d6
`define GTF_CHANNEL__RXLPM_OS_CFG1_SZ 16

`define GTF_CHANNEL__RXOSCALRESET_TIME    32'h000000d7
`define GTF_CHANNEL__RXOSCALRESET_TIME_SZ 5

`define GTF_CHANNEL__RXOUT_DIV    32'h000000d8
`define GTF_CHANNEL__RXOUT_DIV_SZ 6

`define GTF_CHANNEL__RXPCSRESET_TIME    32'h000000d9
`define GTF_CHANNEL__RXPCSRESET_TIME_SZ 5

`define GTF_CHANNEL__RXPHBEACON_CFG    32'h000000da
`define GTF_CHANNEL__RXPHBEACON_CFG_SZ 16

`define GTF_CHANNEL__RXPHBEACON_RAW_CFG    32'h000000db
`define GTF_CHANNEL__RXPHBEACON_RAW_CFG_SZ 16

`define GTF_CHANNEL__RXPHDLY_CFG    32'h000000dc
`define GTF_CHANNEL__RXPHDLY_CFG_SZ 16

`define GTF_CHANNEL__RXPHSAMP_CFG    32'h000000dd
`define GTF_CHANNEL__RXPHSAMP_CFG_SZ 16

`define GTF_CHANNEL__RXPHSAMP_RAW_CFG    32'h000000de
`define GTF_CHANNEL__RXPHSAMP_RAW_CFG_SZ 16

`define GTF_CHANNEL__RXPHSLIP_CFG    32'h000000df
`define GTF_CHANNEL__RXPHSLIP_CFG_SZ 16

`define GTF_CHANNEL__RXPHSLIP_RAW_CFG    32'h000000e0
`define GTF_CHANNEL__RXPHSLIP_RAW_CFG_SZ 16

`define GTF_CHANNEL__RXPH_MONITOR_SEL    32'h000000e1
`define GTF_CHANNEL__RXPH_MONITOR_SEL_SZ 5

`define GTF_CHANNEL__RXPI_CFG0    32'h000000e2
`define GTF_CHANNEL__RXPI_CFG0_SZ 16

`define GTF_CHANNEL__RXPI_CFG1    32'h000000e3
`define GTF_CHANNEL__RXPI_CFG1_SZ 16

`define GTF_CHANNEL__RXPMACLK_SEL    32'h000000e4
`define GTF_CHANNEL__RXPMACLK_SEL_SZ 64

`define GTF_CHANNEL__RXPMARESET_TIME    32'h000000e5
`define GTF_CHANNEL__RXPMARESET_TIME_SZ 5

`define GTF_CHANNEL__RXPRBS_ERR_LOOPBACK    32'h000000e6
`define GTF_CHANNEL__RXPRBS_ERR_LOOPBACK_SZ 1

`define GTF_CHANNEL__RXPRBS_LINKACQ_CNT    32'h000000e7
`define GTF_CHANNEL__RXPRBS_LINKACQ_CNT_SZ 8

`define GTF_CHANNEL__RXREFCLKDIV2_SEL    32'h000000e8
`define GTF_CHANNEL__RXREFCLKDIV2_SEL_SZ 1

`define GTF_CHANNEL__RXSLIDE_AUTO_WAIT    32'h000000e9
`define GTF_CHANNEL__RXSLIDE_AUTO_WAIT_SZ 4

`define GTF_CHANNEL__RXSLIDE_MODE    32'h000000ea
`define GTF_CHANNEL__RXSLIDE_MODE_SZ 32

`define GTF_CHANNEL__RXSYNC_MULTILANE    32'h000000eb
`define GTF_CHANNEL__RXSYNC_MULTILANE_SZ 1

`define GTF_CHANNEL__RXSYNC_OVRD    32'h000000ec
`define GTF_CHANNEL__RXSYNC_OVRD_SZ 1

`define GTF_CHANNEL__RXSYNC_SKIP_DA    32'h000000ed
`define GTF_CHANNEL__RXSYNC_SKIP_DA_SZ 1

`define GTF_CHANNEL__RX_AFE_CM_EN    32'h000000ee
`define GTF_CHANNEL__RX_AFE_CM_EN_SZ 1

`define GTF_CHANNEL__RX_BIAS_CFG0    32'h000000ef
`define GTF_CHANNEL__RX_BIAS_CFG0_SZ 16

`define GTF_CHANNEL__RX_CAPFF_SARC_ENB    32'h000000f0
`define GTF_CHANNEL__RX_CAPFF_SARC_ENB_SZ 1

`define GTF_CHANNEL__RX_CLK25_DIV    32'h000000f1
`define GTF_CHANNEL__RX_CLK25_DIV_SZ 6

`define GTF_CHANNEL__RX_CLKMUX_EN    32'h000000f2
`define GTF_CHANNEL__RX_CLKMUX_EN_SZ 1

`define GTF_CHANNEL__RX_CLK_SLIP_OVRD    32'h000000f3
`define GTF_CHANNEL__RX_CLK_SLIP_OVRD_SZ 5

`define GTF_CHANNEL__RX_CM_BUF_CFG    32'h000000f4
`define GTF_CHANNEL__RX_CM_BUF_CFG_SZ 4

`define GTF_CHANNEL__RX_CM_BUF_PD    32'h000000f5
`define GTF_CHANNEL__RX_CM_BUF_PD_SZ 1

`define GTF_CHANNEL__RX_CM_SEL    32'h000000f6
`define GTF_CHANNEL__RX_CM_SEL_SZ 2

`define GTF_CHANNEL__RX_CM_TRIM    32'h000000f7
`define GTF_CHANNEL__RX_CM_TRIM_SZ 4

`define GTF_CHANNEL__RX_CTLE_PWR_SAVING    32'h000000f8
`define GTF_CHANNEL__RX_CTLE_PWR_SAVING_SZ 1

`define GTF_CHANNEL__RX_CTLE_RES_CTRL    32'h000000f9
`define GTF_CHANNEL__RX_CTLE_RES_CTRL_SZ 4

`define GTF_CHANNEL__RX_DATA_WIDTH    32'h000000fa
`define GTF_CHANNEL__RX_DATA_WIDTH_SZ 8

`define GTF_CHANNEL__RX_DDI_SEL    32'h000000fb
`define GTF_CHANNEL__RX_DDI_SEL_SZ 6

`define GTF_CHANNEL__RX_DEGEN_CTRL    32'h000000fc
`define GTF_CHANNEL__RX_DEGEN_CTRL_SZ 3

`define GTF_CHANNEL__RX_DFELPM_CFG0    32'h000000fd
`define GTF_CHANNEL__RX_DFELPM_CFG0_SZ 4

`define GTF_CHANNEL__RX_DFELPM_CFG1    32'h000000fe
`define GTF_CHANNEL__RX_DFELPM_CFG1_SZ 1

`define GTF_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN    32'h000000ff
`define GTF_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN_SZ 1

`define GTF_CHANNEL__RX_DFE_AGC_CFG1    32'h00000100
`define GTF_CHANNEL__RX_DFE_AGC_CFG1_SZ 3

`define GTF_CHANNEL__RX_DFE_KL_LPM_KH_CFG0    32'h00000101
`define GTF_CHANNEL__RX_DFE_KL_LPM_KH_CFG0_SZ 2

`define GTF_CHANNEL__RX_DFE_KL_LPM_KH_CFG1    32'h00000102
`define GTF_CHANNEL__RX_DFE_KL_LPM_KH_CFG1_SZ 3

`define GTF_CHANNEL__RX_DFE_KL_LPM_KL_CFG0    32'h00000103
`define GTF_CHANNEL__RX_DFE_KL_LPM_KL_CFG0_SZ 2

`define GTF_CHANNEL__RX_DFE_KL_LPM_KL_CFG1    32'h00000104
`define GTF_CHANNEL__RX_DFE_KL_LPM_KL_CFG1_SZ 3

`define GTF_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE    32'h00000105
`define GTF_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE_SZ 1

`define GTF_CHANNEL__RX_DISPERR_SEQ_MATCH    32'h00000106
`define GTF_CHANNEL__RX_DISPERR_SEQ_MATCH_SZ 40

`define GTF_CHANNEL__RX_DIVRESET_TIME    32'h00000107
`define GTF_CHANNEL__RX_DIVRESET_TIME_SZ 5

`define GTF_CHANNEL__RX_EN_CTLE_RCAL_B    32'h00000108
`define GTF_CHANNEL__RX_EN_CTLE_RCAL_B_SZ 1

`define GTF_CHANNEL__RX_EN_SUM_RCAL_B    32'h00000109
`define GTF_CHANNEL__RX_EN_SUM_RCAL_B_SZ 1

`define GTF_CHANNEL__RX_EYESCAN_VS_CODE    32'h0000010a
`define GTF_CHANNEL__RX_EYESCAN_VS_CODE_SZ 7

`define GTF_CHANNEL__RX_EYESCAN_VS_NEG_DIR    32'h0000010b
`define GTF_CHANNEL__RX_EYESCAN_VS_NEG_DIR_SZ 1

`define GTF_CHANNEL__RX_EYESCAN_VS_RANGE    32'h0000010c
`define GTF_CHANNEL__RX_EYESCAN_VS_RANGE_SZ 2

`define GTF_CHANNEL__RX_EYESCAN_VS_UT_SIGN    32'h0000010d
`define GTF_CHANNEL__RX_EYESCAN_VS_UT_SIGN_SZ 1

`define GTF_CHANNEL__RX_I2V_FILTER_EN    32'h0000010e
`define GTF_CHANNEL__RX_I2V_FILTER_EN_SZ 1

`define GTF_CHANNEL__RX_INT_DATAWIDTH    32'h0000010f
`define GTF_CHANNEL__RX_INT_DATAWIDTH_SZ 2

`define GTF_CHANNEL__RX_PMA_POWER_SAVE    32'h00000110
`define GTF_CHANNEL__RX_PMA_POWER_SAVE_SZ 1

`define GTF_CHANNEL__RX_PMA_RSV0    32'h00000111
`define GTF_CHANNEL__RX_PMA_RSV0_SZ 16

`define GTF_CHANNEL__RX_PROGDIV_CFG    32'h00000112
`define GTF_CHANNEL__RX_PROGDIV_CFG_SZ 64

`define GTF_CHANNEL__RX_PROGDIV_RATE    32'h00000113
`define GTF_CHANNEL__RX_PROGDIV_RATE_SZ 16

`define GTF_CHANNEL__RX_RESLOAD_CTRL    32'h00000114
`define GTF_CHANNEL__RX_RESLOAD_CTRL_SZ 4

`define GTF_CHANNEL__RX_RESLOAD_OVRD    32'h00000115
`define GTF_CHANNEL__RX_RESLOAD_OVRD_SZ 1

`define GTF_CHANNEL__RX_SAMPLE_PERIOD    32'h00000116
`define GTF_CHANNEL__RX_SAMPLE_PERIOD_SZ 3

`define GTF_CHANNEL__RX_SIG_VALID_DLY    32'h00000117
`define GTF_CHANNEL__RX_SIG_VALID_DLY_SZ 6

`define GTF_CHANNEL__RX_SUM_DEGEN_AVTT_OVERITE    32'h00000118
`define GTF_CHANNEL__RX_SUM_DEGEN_AVTT_OVERITE_SZ 1

`define GTF_CHANNEL__RX_SUM_DFETAPREP_EN    32'h00000119
`define GTF_CHANNEL__RX_SUM_DFETAPREP_EN_SZ 1

`define GTF_CHANNEL__RX_SUM_IREF_TUNE    32'h0000011a
`define GTF_CHANNEL__RX_SUM_IREF_TUNE_SZ 4

`define GTF_CHANNEL__RX_SUM_PWR_SAVING    32'h0000011b
`define GTF_CHANNEL__RX_SUM_PWR_SAVING_SZ 1

`define GTF_CHANNEL__RX_SUM_RES_CTRL    32'h0000011c
`define GTF_CHANNEL__RX_SUM_RES_CTRL_SZ 4

`define GTF_CHANNEL__RX_SUM_VCMTUNE    32'h0000011d
`define GTF_CHANNEL__RX_SUM_VCMTUNE_SZ 4

`define GTF_CHANNEL__RX_SUM_VCM_BIAS_TUNE_EN    32'h0000011e
`define GTF_CHANNEL__RX_SUM_VCM_BIAS_TUNE_EN_SZ 1

`define GTF_CHANNEL__RX_SUM_VCM_OVWR    32'h0000011f
`define GTF_CHANNEL__RX_SUM_VCM_OVWR_SZ 1

`define GTF_CHANNEL__RX_SUM_VREF_TUNE    32'h00000120
`define GTF_CHANNEL__RX_SUM_VREF_TUNE_SZ 3

`define GTF_CHANNEL__RX_TUNE_AFE_OS    32'h00000121
`define GTF_CHANNEL__RX_TUNE_AFE_OS_SZ 2

`define GTF_CHANNEL__RX_VREG_CTRL    32'h00000122
`define GTF_CHANNEL__RX_VREG_CTRL_SZ 3

`define GTF_CHANNEL__RX_VREG_PDB    32'h00000123
`define GTF_CHANNEL__RX_VREG_PDB_SZ 1

`define GTF_CHANNEL__RX_WIDEMODE_CDR    32'h00000124
`define GTF_CHANNEL__RX_WIDEMODE_CDR_SZ 2

`define GTF_CHANNEL__RX_WIDEMODE_CDR_GEN3    32'h00000125
`define GTF_CHANNEL__RX_WIDEMODE_CDR_GEN3_SZ 2

`define GTF_CHANNEL__RX_WIDEMODE_CDR_GEN4    32'h00000126
`define GTF_CHANNEL__RX_WIDEMODE_CDR_GEN4_SZ 2

`define GTF_CHANNEL__RX_XCLK_SEL    32'h00000127
`define GTF_CHANNEL__RX_XCLK_SEL_SZ 40

`define GTF_CHANNEL__RX_XMODE_SEL    32'h00000128
`define GTF_CHANNEL__RX_XMODE_SEL_SZ 1

`define GTF_CHANNEL__SAMPLE_CLK_PHASE    32'h00000129
`define GTF_CHANNEL__SAMPLE_CLK_PHASE_SZ 1

`define GTF_CHANNEL__SATA_CPLL_CFG    32'h0000012a
`define GTF_CHANNEL__SATA_CPLL_CFG_SZ 88

`define GTF_CHANNEL__SIM_MODE    32'h0000012b
`define GTF_CHANNEL__SIM_MODE_SZ 48

`define GTF_CHANNEL__SIM_RESET_SPEEDUP    32'h0000012c
`define GTF_CHANNEL__SIM_RESET_SPEEDUP_SZ 40

`define GTF_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL    32'h0000012d
`define GTF_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTF_CHANNEL__SRSTMODE    32'h0000012e
`define GTF_CHANNEL__SRSTMODE_SZ 1

`define GTF_CHANNEL__TAPDLY_SET_TX    32'h0000012f
`define GTF_CHANNEL__TAPDLY_SET_TX_SZ 2

`define GTF_CHANNEL__TCO_NEW_CFG0    32'h00000130
`define GTF_CHANNEL__TCO_NEW_CFG0_SZ 16

`define GTF_CHANNEL__TCO_NEW_CFG1    32'h00000131
`define GTF_CHANNEL__TCO_NEW_CFG1_SZ 16

`define GTF_CHANNEL__TCO_NEW_CFG2    32'h00000132
`define GTF_CHANNEL__TCO_NEW_CFG2_SZ 16

`define GTF_CHANNEL__TCO_NEW_CFG3    32'h00000133
`define GTF_CHANNEL__TCO_NEW_CFG3_SZ 16

`define GTF_CHANNEL__TCO_RSVD1    32'h00000134
`define GTF_CHANNEL__TCO_RSVD1_SZ 16

`define GTF_CHANNEL__TCO_RSVD2    32'h00000135
`define GTF_CHANNEL__TCO_RSVD2_SZ 16

`define GTF_CHANNEL__TERM_RCAL_CFG    32'h00000136
`define GTF_CHANNEL__TERM_RCAL_CFG_SZ 15

`define GTF_CHANNEL__TERM_RCAL_OVRD    32'h00000137
`define GTF_CHANNEL__TERM_RCAL_OVRD_SZ 3

`define GTF_CHANNEL__TRANS_TIME_RATE    32'h00000138
`define GTF_CHANNEL__TRANS_TIME_RATE_SZ 8

`define GTF_CHANNEL__TST_RSV0    32'h00000139
`define GTF_CHANNEL__TST_RSV0_SZ 8

`define GTF_CHANNEL__TST_RSV1    32'h0000013a
`define GTF_CHANNEL__TST_RSV1_SZ 8

`define GTF_CHANNEL__TXBUF_EN    32'h0000013b
`define GTF_CHANNEL__TXBUF_EN_SZ 40

`define GTF_CHANNEL__TXDLY_CFG    32'h0000013c
`define GTF_CHANNEL__TXDLY_CFG_SZ 16

`define GTF_CHANNEL__TXDLY_LCFG    32'h0000013d
`define GTF_CHANNEL__TXDLY_LCFG_SZ 16

`define GTF_CHANNEL__TXDRV_FREQBAND    32'h0000013e
`define GTF_CHANNEL__TXDRV_FREQBAND_SZ 2

`define GTF_CHANNEL__TXFE_CFG0    32'h0000013f
`define GTF_CHANNEL__TXFE_CFG0_SZ 16

`define GTF_CHANNEL__TXFE_CFG1    32'h00000140
`define GTF_CHANNEL__TXFE_CFG1_SZ 16

`define GTF_CHANNEL__TXFE_CFG2    32'h00000141
`define GTF_CHANNEL__TXFE_CFG2_SZ 16

`define GTF_CHANNEL__TXFE_CFG3    32'h00000142
`define GTF_CHANNEL__TXFE_CFG3_SZ 16

`define GTF_CHANNEL__TXFIFO_ADDR_CFG    32'h00000143
`define GTF_CHANNEL__TXFIFO_ADDR_CFG_SZ 32

`define GTF_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR    32'h00000144
`define GTF_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR_SZ 3

`define GTF_CHANNEL__TXOUT_DIV    32'h00000145
`define GTF_CHANNEL__TXOUT_DIV_SZ 6

`define GTF_CHANNEL__TXPCSRESET_TIME    32'h00000146
`define GTF_CHANNEL__TXPCSRESET_TIME_SZ 5

`define GTF_CHANNEL__TXPHDLY_CFG0    32'h00000147
`define GTF_CHANNEL__TXPHDLY_CFG0_SZ 16

`define GTF_CHANNEL__TXPHDLY_CFG1    32'h00000148
`define GTF_CHANNEL__TXPHDLY_CFG1_SZ 16

`define GTF_CHANNEL__TXPH_CFG    32'h00000149
`define GTF_CHANNEL__TXPH_CFG_SZ 16

`define GTF_CHANNEL__TXPH_CFG2    32'h0000014a
`define GTF_CHANNEL__TXPH_CFG2_SZ 16

`define GTF_CHANNEL__TXPH_MONITOR_SEL    32'h0000014b
`define GTF_CHANNEL__TXPH_MONITOR_SEL_SZ 5

`define GTF_CHANNEL__TXPI_CFG0    32'h0000014c
`define GTF_CHANNEL__TXPI_CFG0_SZ 16

`define GTF_CHANNEL__TXPI_CFG1    32'h0000014d
`define GTF_CHANNEL__TXPI_CFG1_SZ 16

`define GTF_CHANNEL__TXPI_GRAY_SEL    32'h0000014e
`define GTF_CHANNEL__TXPI_GRAY_SEL_SZ 1

`define GTF_CHANNEL__TXPI_INVSTROBE_SEL    32'h0000014f
`define GTF_CHANNEL__TXPI_INVSTROBE_SEL_SZ 1

`define GTF_CHANNEL__TXPI_PPM    32'h00000150
`define GTF_CHANNEL__TXPI_PPM_SZ 1

`define GTF_CHANNEL__TXPI_PPM_CFG    32'h00000151
`define GTF_CHANNEL__TXPI_PPM_CFG_SZ 8

`define GTF_CHANNEL__TXPI_SYNFREQ_PPM    32'h00000152
`define GTF_CHANNEL__TXPI_SYNFREQ_PPM_SZ 3

`define GTF_CHANNEL__TXPMARESET_TIME    32'h00000153
`define GTF_CHANNEL__TXPMARESET_TIME_SZ 5

`define GTF_CHANNEL__TXREFCLKDIV2_SEL    32'h00000154
`define GTF_CHANNEL__TXREFCLKDIV2_SEL_SZ 1

`define GTF_CHANNEL__TXSWBST_BST    32'h00000155
`define GTF_CHANNEL__TXSWBST_BST_SZ 2

`define GTF_CHANNEL__TXSWBST_EN    32'h00000156
`define GTF_CHANNEL__TXSWBST_EN_SZ 1

`define GTF_CHANNEL__TXSWBST_MAG    32'h00000157
`define GTF_CHANNEL__TXSWBST_MAG_SZ 3

`define GTF_CHANNEL__TXSYNC_MULTILANE    32'h00000158
`define GTF_CHANNEL__TXSYNC_MULTILANE_SZ 1

`define GTF_CHANNEL__TXSYNC_OVRD    32'h00000159
`define GTF_CHANNEL__TXSYNC_OVRD_SZ 1

`define GTF_CHANNEL__TXSYNC_SKIP_DA    32'h0000015a
`define GTF_CHANNEL__TXSYNC_SKIP_DA_SZ 1

`define GTF_CHANNEL__TX_CLK25_DIV    32'h0000015b
`define GTF_CHANNEL__TX_CLK25_DIV_SZ 6

`define GTF_CHANNEL__TX_CLKMUX_EN    32'h0000015c
`define GTF_CHANNEL__TX_CLKMUX_EN_SZ 1

`define GTF_CHANNEL__TX_DATA_WIDTH    32'h0000015d
`define GTF_CHANNEL__TX_DATA_WIDTH_SZ 8

`define GTF_CHANNEL__TX_DCC_LOOP_RST_CFG    32'h0000015e
`define GTF_CHANNEL__TX_DCC_LOOP_RST_CFG_SZ 16

`define GTF_CHANNEL__TX_DIVRESET_TIME    32'h0000015f
`define GTF_CHANNEL__TX_DIVRESET_TIME_SZ 5

`define GTF_CHANNEL__TX_EIDLE_ASSERT_DELAY    32'h00000160
`define GTF_CHANNEL__TX_EIDLE_ASSERT_DELAY_SZ 3

`define GTF_CHANNEL__TX_EIDLE_DEASSERT_DELAY    32'h00000161
`define GTF_CHANNEL__TX_EIDLE_DEASSERT_DELAY_SZ 3

`define GTF_CHANNEL__TX_FABINT_USRCLK_FLOP    32'h00000162
`define GTF_CHANNEL__TX_FABINT_USRCLK_FLOP_SZ 1

`define GTF_CHANNEL__TX_FIFO_BYP_EN    32'h00000163
`define GTF_CHANNEL__TX_FIFO_BYP_EN_SZ 1

`define GTF_CHANNEL__TX_IDLE_DATA_ZERO    32'h00000164
`define GTF_CHANNEL__TX_IDLE_DATA_ZERO_SZ 1

`define GTF_CHANNEL__TX_INT_DATAWIDTH    32'h00000165
`define GTF_CHANNEL__TX_INT_DATAWIDTH_SZ 2

`define GTF_CHANNEL__TX_LOOPBACK_DRIVE_HIZ    32'h00000166
`define GTF_CHANNEL__TX_LOOPBACK_DRIVE_HIZ_SZ 40

`define GTF_CHANNEL__TX_MAINCURSOR_SEL    32'h00000167
`define GTF_CHANNEL__TX_MAINCURSOR_SEL_SZ 1

`define GTF_CHANNEL__TX_PHICAL_CFG0    32'h00000168
`define GTF_CHANNEL__TX_PHICAL_CFG0_SZ 16

`define GTF_CHANNEL__TX_PHICAL_CFG1    32'h00000169
`define GTF_CHANNEL__TX_PHICAL_CFG1_SZ 16

`define GTF_CHANNEL__TX_PI_BIASSET    32'h0000016a
`define GTF_CHANNEL__TX_PI_BIASSET_SZ 2

`define GTF_CHANNEL__TX_PMADATA_OPT    32'h0000016b
`define GTF_CHANNEL__TX_PMADATA_OPT_SZ 1

`define GTF_CHANNEL__TX_PMA_POWER_SAVE    32'h0000016c
`define GTF_CHANNEL__TX_PMA_POWER_SAVE_SZ 1

`define GTF_CHANNEL__TX_PMA_RSV0    32'h0000016d
`define GTF_CHANNEL__TX_PMA_RSV0_SZ 16

`define GTF_CHANNEL__TX_PMA_RSV1    32'h0000016e
`define GTF_CHANNEL__TX_PMA_RSV1_SZ 16

`define GTF_CHANNEL__TX_PROGCLK_SEL    32'h0000016f
`define GTF_CHANNEL__TX_PROGCLK_SEL_SZ 48

`define GTF_CHANNEL__TX_PROGDIV_CFG    32'h00000170
`define GTF_CHANNEL__TX_PROGDIV_CFG_SZ 64

`define GTF_CHANNEL__TX_PROGDIV_RATE    32'h00000171
`define GTF_CHANNEL__TX_PROGDIV_RATE_SZ 16

`define GTF_CHANNEL__TX_SAMPLE_PERIOD    32'h00000172
`define GTF_CHANNEL__TX_SAMPLE_PERIOD_SZ 3

`define GTF_CHANNEL__TX_SW_MEAS    32'h00000173
`define GTF_CHANNEL__TX_SW_MEAS_SZ 2

`define GTF_CHANNEL__TX_VREG_CTRL    32'h00000174
`define GTF_CHANNEL__TX_VREG_CTRL_SZ 3

`define GTF_CHANNEL__TX_VREG_PDB    32'h00000175
`define GTF_CHANNEL__TX_VREG_PDB_SZ 1

`define GTF_CHANNEL__TX_VREG_VREFSEL    32'h00000176
`define GTF_CHANNEL__TX_VREG_VREFSEL_SZ 2

`define GTF_CHANNEL__TX_XCLK_SEL    32'h00000177
`define GTF_CHANNEL__TX_XCLK_SEL_SZ 40

`define GTF_CHANNEL__USE_PCS_CLK_PHASE_SEL    32'h00000178
`define GTF_CHANNEL__USE_PCS_CLK_PHASE_SEL_SZ 1

`define GTF_CHANNEL__USE_RAW_ELEC    32'h00000179
`define GTF_CHANNEL__USE_RAW_ELEC_SZ 1

`define GTF_CHANNEL__Y_ALL_MODE    32'h0000017a
`define GTF_CHANNEL__Y_ALL_MODE_SZ 1

`endif  // B_GTF_CHANNEL_DEFINES_VH