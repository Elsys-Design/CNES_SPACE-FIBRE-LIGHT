`include "B_RFADC_defines.vh"

reg [`RFADC_DATA_SZ-1:0] ATTR [0:`RFADC_ADDR_N-1];
reg [`RFADC__LD_DEVICE_SZ-1:0] LD_DEVICE_REG = LD_DEVICE;
reg [`RFADC__OPT_ANALOG_SZ-1:0] OPT_ANALOG_REG = OPT_ANALOG;
reg [`RFADC__OPT_CLK_DIST_SZ-1:0] OPT_CLK_DIST_REG = OPT_CLK_DIST;
reg [`RFADC__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`RFADC__XPA_ACTIVE_DUTYCYCLE_SZ-1:0] XPA_ACTIVE_DUTYCYCLE_REG = XPA_ACTIVE_DUTYCYCLE;
reg [`RFADC__XPA_CFG0_SZ-1:0] XPA_CFG0_REG = XPA_CFG0;
reg [`RFADC__XPA_CFG1_SZ-1:0] XPA_CFG1_REG = XPA_CFG1;
reg [`RFADC__XPA_CFG2_SZ-1:0] XPA_CFG2_REG = XPA_CFG2;
reg [`RFADC__XPA_NUM_ADCS_SZ:1] XPA_NUM_ADCS_REG = XPA_NUM_ADCS;
reg [`RFADC__XPA_NUM_DDCS_SZ-1:0] XPA_NUM_DDCS_REG = XPA_NUM_DDCS;
reg [`RFADC__XPA_PLL_USED_SZ:1] XPA_PLL_USED_REG = XPA_PLL_USED;
reg [`RFADC__XPA_SAMPLE_RATE_MSPS_SZ-1:0] XPA_SAMPLE_RATE_MSPS_REG = XPA_SAMPLE_RATE_MSPS;

initial begin
  ATTR[`RFADC__LD_DEVICE] = LD_DEVICE;
  ATTR[`RFADC__OPT_ANALOG] = OPT_ANALOG;
  ATTR[`RFADC__OPT_CLK_DIST] = OPT_CLK_DIST;
  ATTR[`RFADC__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`RFADC__XPA_ACTIVE_DUTYCYCLE] = XPA_ACTIVE_DUTYCYCLE;
  ATTR[`RFADC__XPA_CFG0] = XPA_CFG0;
  ATTR[`RFADC__XPA_CFG1] = XPA_CFG1;
  ATTR[`RFADC__XPA_CFG2] = XPA_CFG2;
  ATTR[`RFADC__XPA_NUM_ADCS] = XPA_NUM_ADCS;
  ATTR[`RFADC__XPA_NUM_DDCS] = XPA_NUM_DDCS;
  ATTR[`RFADC__XPA_PLL_USED] = XPA_PLL_USED;
  ATTR[`RFADC__XPA_SAMPLE_RATE_MSPS] = XPA_SAMPLE_RATE_MSPS;
end

always @(trig_attr) begin
  LD_DEVICE_REG = ATTR[`RFADC__LD_DEVICE];
  OPT_ANALOG_REG = ATTR[`RFADC__OPT_ANALOG];
  OPT_CLK_DIST_REG = ATTR[`RFADC__OPT_CLK_DIST];
  SIM_DEVICE_REG = ATTR[`RFADC__SIM_DEVICE];
  XPA_ACTIVE_DUTYCYCLE_REG = ATTR[`RFADC__XPA_ACTIVE_DUTYCYCLE];
  XPA_CFG0_REG = ATTR[`RFADC__XPA_CFG0];
  XPA_CFG1_REG = ATTR[`RFADC__XPA_CFG1];
  XPA_CFG2_REG = ATTR[`RFADC__XPA_CFG2];
  XPA_NUM_ADCS_REG = ATTR[`RFADC__XPA_NUM_ADCS];
  XPA_NUM_DDCS_REG = ATTR[`RFADC__XPA_NUM_DDCS];
  XPA_PLL_USED_REG = ATTR[`RFADC__XPA_PLL_USED];
  XPA_SAMPLE_RATE_MSPS_REG = ATTR[`RFADC__XPA_SAMPLE_RATE_MSPS];
end

// procedures to override, read attribute values

task write_attr;
  input  [`RFADC_ADDR_SZ-1:0] addr;
  input  [`RFADC_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`RFADC_DATA_SZ-1:0] read_attr;
  input  [`RFADC_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
