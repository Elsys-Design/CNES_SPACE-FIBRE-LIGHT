-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 16/07/2025
--
-- Description : This module inserts control words into the data flow
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_lane_ctrl_word_insert is
  port (
    RST_N                                : in  std_logic;                                   --! Global reset Active Low
    CLK                                  : in  std_logic;                                   --! Clock generated by HSSL IP
    -- Data-Link interface
    RD_DATA_EN_PLCWI                     : out std_logic;                                   --! Read command to receive data from the Data-Link layer
    RD_DATA_VALID_DL                     : in  std_logic;                                   --! Data valid flag from the Data-Link layer
    CAPABILITY_DL                        : in  std_logic_vector(7 downto 0);                --! Capability field from the Data-Link layer
    DATA_TX_DL                           : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data received from the Data-Link layer
    VALID_K_CHARAC_DL                    : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicating which bytes are K characters from the Data-Link layer
    NO_DATA_DL                           : in  std_logic;                                   --! Flag enabling IDLE word insertion when no data is available from the Data-Link layer
    -- ppl_64_skip_insertion (PLSI) interface
    WAIT_SEND_DATA_PLSI                  : in  std_logic;                                   --! Flag indicating that skip_insertion is sending a SKIP control word
    NEW_DATA_PLCWI                       : out std_logic;                                   --! New data available for skip_insertion
    DATA_TX_PLCWI                        : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to be sent to the physical layer
    VALID_K_CHARAC_PLCWI                 : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicating which bytes are K characters
    -- ppl_64_lane_init_fsm (PLIF) interface
    SEND_INIT1_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT1 control word followed by 64 pseudo-random data words
    SEND_INIT2_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT2 control word followed by 64 pseudo-random data words
    SEND_INIT3_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT3 control word followed by 64 pseudo-random data words
    ENABLE_TRANSM_DATA_PLIF              : in  std_logic;                                   --! Flag to enable data transmission
    SEND_32_STANDBY_CTRL_WORDS_PLIF      : in  std_logic;                                   --! Flag to send 32 STANDBY control words
    SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF  : in  std_logic;                                   --! Flag to send 32 LOSS_SIGNAL control words
    STANDBY_SIGNAL_X32_PLCWI             : out std_logic;                                   --! Flag indicating 32 STANDBY control words have been sent
    LOST_SIGNAL_X32_PLCWI                : out std_logic;                                   --! Flag indicating 32 LOSS_SIGNAL control words have been sent
    LOST_CAUSE_PLIF                      : in  std_logic_vector(1 downto 0);                --! Indicates the reason for LOST_SIGNAL
    -- MIB interface
    STANDBY_REASON_MIB                   : in  std_logic_vector(7 downto 0)                 --! Standby reason from MIB
  );
end ppl_64_lane_ctrl_word_insert;

architecture rtl of ppl_64_lane_ctrl_word_insert is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------

signal prbs_counter      : unsigned(31 downto 0);
signal send_stdby_cnt    : unsigned(5 downto 0);
signal send_loss_sig_cnt : unsigned(5 downto 0);
signal no_data_dl_r      : std_logic;

begin

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_send_data
--! Inserts conrtol words into the data flow 
---------------------------------------------------------
  p_send_data : process(CLK, RST_N)
  begin
    if RST_N = '0' then
      RD_DATA_EN_PLCWI               <= '0';
      NEW_DATA_PLCWI                 <= '0';
      DATA_TX_PLCWI                  <= (others => '0');
      VALID_K_CHARAC_PLCWI           <= (others => '0');
      prbs_counter                   <= (others => '0');
      send_stdby_cnt                 <= (others => '0');
      STANDBY_SIGNAL_X32_PLCWI       <= '0';
      send_loss_sig_cnt              <= (others => '0');
      LOST_SIGNAL_X32_PLCWI          <= '0';
      no_data_dl_r                   <= '0';
    elsif rising_edge(CLK) then
      no_data_dl_r                   <= NO_DATA_DL;
      RD_DATA_EN_PLCWI               <= '0';
      STANDBY_SIGNAL_X32_PLCWI       <= '0';
      LOST_SIGNAL_X32_PLCWI          <= '0';

      --------------------------------------
      --          INIT Control Word        --
      --------------------------------------
      if SEND_INIT1_CTRL_WORD_PLIF = '1' or SEND_INIT2_CTRL_WORD_PLIF = '1' or SEND_INIT3_CTRL_WORD_PLIF = '1' then
        if prbs_counter < C_PRBS_COUNTER_64-1 then
          -- Send PRBS
          prbs_counter          <= prbs_counter + 2;  -- 2 PRBS words
          NEW_DATA_PLCWI        <= '1';
          DATA_TX_PLCWI         <= std_logic_vector(prbs_counter + 1) & std_logic_vector(prbs_counter);
          VALID_K_CHARAC_PLCWI  <= x"00";
        elsif prbs_counter = C_PRBS_COUNTER_64-1 then
          -- Insert INIT word on word 2
          NEW_DATA_PLCWI        <= '1';
          VALID_K_CHARAC_PLCWI  <= x"10";
          prbs_counter          <= (others => '0');
          if SEND_INIT1_CTRL_WORD_PLIF = '1' then
            -- Send INIT1 control word
            DATA_TX_PLCWI <= C_INIT1_WORD & std_logic_vector(prbs_counter);
          elsif SEND_INIT2_CTRL_WORD_PLIF = '1' then
            -- Send INIT2 control word
            DATA_TX_PLCWI <= C_INIT2_WORD & std_logic_vector(prbs_counter);
          elsif SEND_INIT3_CTRL_WORD_PLIF = '1' then
            -- Send INIT3 control word
            DATA_TX_PLCWI <= CAPABILITY_DL & C_INIT3_WORD & std_logic_vector(prbs_counter);
          end if;
        elsif prbs_counter = C_PRBS_COUNTER_64 then
          -- Insert INIT word on word 1
          NEW_DATA_PLCWI        <= '1';
          VALID_K_CHARAC_PLCWI  <= x"01";
          prbs_counter          <= to_unsigned(1, prbs_counter'length);
          if SEND_INIT1_CTRL_WORD_PLIF = '1' then
            -- Send INIT1 control word
            DATA_TX_PLCWI       <= x"00000000" & C_INIT1_WORD;
          elsif SEND_INIT2_CTRL_WORD_PLIF = '1' then
            -- Send INIT2 control word
            DATA_TX_PLCWI       <= x"00000000" & C_INIT2_WORD;
          elsif SEND_INIT3_CTRL_WORD_PLIF = '1' then
            -- Send INIT3 control word
            DATA_TX_PLCWI       <= x"00000000" & CAPABILITY_DL & C_INIT3_WORD;
          end if;
        end if;

      --------------------------------------
      --       Active State: Data TX      --
      --------------------------------------
      elsif ENABLE_TRANSM_DATA_PLIF = '1' then
        -- When lane_init_fsm is in ACTIVE_ST
        NEW_DATA_PLCWI <= '1';
        if ((no_data_dl_r = '0' and NO_DATA_DL = '1') or NO_DATA_DL = '0') and WAIT_SEND_DATA_PLSI = '0' then
          RD_DATA_EN_PLCWI <= '1';
          if RD_DATA_VALID_DL = '1' then
            DATA_TX_PLCWI        <= DATA_TX_DL;
            VALID_K_CHARAC_PLCWI <= VALID_K_CHARAC_DL;
          else
            DATA_TX_PLCWI        <= C_IDLE_WORD & C_IDLE_WORD;
            VALID_K_CHARAC_PLCWI <= x"11";
          end if;
        elsif ((no_data_dl_r = '0' and NO_DATA_DL = '1') or NO_DATA_DL = '0') and WAIT_SEND_DATA_PLSI = '1' then
          RD_DATA_EN_PLCWI <= '0';
          if RD_DATA_VALID_DL = '1' then
            DATA_TX_PLCWI        <= DATA_TX_DL;
            VALID_K_CHARAC_PLCWI <= VALID_K_CHARAC_DL;
          else
            DATA_TX_PLCWI        <= C_IDLE_WORD & C_IDLE_WORD;
            VALID_K_CHARAC_PLCWI <= x"11";
          end if;
        else
          -- No data available from the Data-Link layer
          RD_DATA_EN_PLCWI       <= '1';
          DATA_TX_PLCWI          <= C_IDLE_WORD & C_IDLE_WORD;
          VALID_K_CHARAC_PLCWI   <= x"11";
        end if;

      --------------------------------------
      --       STANDBY Control Word       --
      --------------------------------------
      elsif SEND_32_STANDBY_CTRL_WORDS_PLIF = '1' then
        -- When lane_init_fsm is in PREPARE_STANDBY_ST
        if send_stdby_cnt >= C_X32_SIGNAL then
          -- 32 STANDBY control words have been sent
          STANDBY_SIGNAL_X32_PLCWI <= '1';
          send_stdby_cnt           <= (others => '0');
        else
          STANDBY_SIGNAL_X32_PLCWI <= '0';
          send_stdby_cnt           <= send_stdby_cnt + 2;
          NEW_DATA_PLCWI           <= '1';
          DATA_TX_PLCWI            <= STANDBY_REASON_MIB & C_STANDBY_WORD & STANDBY_REASON_MIB & C_STANDBY_WORD;
          VALID_K_CHARAC_PLCWI     <= x"11";
        end if;

      --------------------------------------
      --     LOSS SIGNAL Control Word     --
      --------------------------------------
      elsif SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF = '1' then
        -- When lane_init_fsm is in LOSS_OF_SIGNAL_ST
        if send_loss_sig_cnt >= C_X32_SIGNAL then
          -- 32 LOSS_SIGNAL control words have been sent
          LOST_SIGNAL_X32_PLCWI <= '1';
          send_loss_sig_cnt     <= (others => '0');
        else
          LOST_SIGNAL_X32_PLCWI <= '0';
          send_loss_sig_cnt     <= send_loss_sig_cnt + 2;
          NEW_DATA_PLCWI        <= '1';
          DATA_TX_PLCWI         <= "000000" & LOST_CAUSE_PLIF & C_LOST_SIG_WORD & "000000" & LOST_CAUSE_PLIF & C_LOST_SIG_WORD;
          VALID_K_CHARAC_PLCWI  <= x"11";
        end if;

      else
        NEW_DATA_PLCWI        <= '0';
        DATA_TX_PLCWI         <= (others => '0');
        VALID_K_CHARAC_PLCWI  <= (others => '0');
        prbs_counter          <= (others => '0');
        send_stdby_cnt        <= (others => '0');
        send_loss_sig_cnt     <= (others => '0');
      end if;
    end if;
  end process p_send_data;

end architecture rtl;
