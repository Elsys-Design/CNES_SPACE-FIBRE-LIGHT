// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_FP_OUTPUT_DEFINES_VH
`else
`define B_DSP_FP_OUTPUT_DEFINES_VH

// Look-up table parameters
//

`define DSP_FP_OUTPUT_ADDR_N  7
`define DSP_FP_OUTPUT_ADDR_SZ 32
`define DSP_FP_OUTPUT_DATA_SZ 64

// Attribute addresses
//

`define DSP_FP_OUTPUT__FPA_PREG    32'h00000000
`define DSP_FP_OUTPUT__FPA_PREG_SZ 32

`define DSP_FP_OUTPUT__FPM_PREG    32'h00000001
`define DSP_FP_OUTPUT__FPM_PREG_SZ 32

`define DSP_FP_OUTPUT__IS_RSTFPA_INVERTED    32'h00000002
`define DSP_FP_OUTPUT__IS_RSTFPA_INVERTED_SZ 1

`define DSP_FP_OUTPUT__IS_RSTFPM_INVERTED    32'h00000003
`define DSP_FP_OUTPUT__IS_RSTFPM_INVERTED_SZ 1

`define DSP_FP_OUTPUT__PCOUTSEL    32'h00000004
`define DSP_FP_OUTPUT__PCOUTSEL_SZ 24

`define DSP_FP_OUTPUT__RESET_MODE    32'h00000005
`define DSP_FP_OUTPUT__RESET_MODE_SZ 40

`define DSP_FP_OUTPUT__USE_MULT    32'h00000006
`define DSP_FP_OUTPUT__USE_MULT_SZ 64

`endif  // B_DSP_FP_OUTPUT_DEFINES_VH