-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation data : 03/07/2024
--
--- Description: This module implements the receive synchronization state machine
----------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;
  
entity ppl_64_rx_sync_fsm is
  port(
    RST_N                            : in  std_logic;                                    --! Global reset. Active low
    CLK                              : in  std_logic;                                    --! Clock generated by GTY IP
    -- Data-link layer interface
    LANE_RESET_DL                    : in  std_logic;                                    --! Lane reset command from Data-Link Layer.
    -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
    DATA_RX_PLRSF                    : out std_logic_vector(C_DATA_WIDTH-1  downto 0);   --! 64-bit data to lane_ctrl_word_detect
    VALID_K_CHARAC_PLRSF             : out std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! 8-bit valid K character flags to lane_ctrl_word_detect
    DATA_RDY_PLRSF                   : out std_logic;                                    --! Data valid flag to lane_ctrl_word_detect
    -- ppl_64_word_alignment (PLWA) interface
    DATA_RX_PLWA                     : in  std_logic_vector(C_DATA_WIDTH-1  downto 0);   --! 64-bit data from ppl_64_word_alignment
    VALID_K_CHARAC_PLWA              : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! 8-bit valid K character flags from ppl_64_word_alignment
    INVALID_CHAR_PLWA                : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Invalid character flags from ppl_64_word_alignment
    DISPARITY_ERR_PLWA               : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Disparity error flags from ppl_64_word_alignment
    RX_WORD_IS_ALIGNED_PLWA          : in  std_logic;                                    --! RX word is aligned from ppl_64_word_alignment
    COMMA_DET_PLWA                   : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Flag indicates that a comma is detected on the word received
    -- PARAMETERS (MIB)
    LANE_RESET                       : in  std_logic                                     --! Asserts or de-asserts LaneReset for the lane
  );
end ppl_64_rx_sync_fsm;

architecture rtl of ppl_64_rx_sync_fsm is
---------------------------------------------------------
----- Type declaration -----
---------------------------------------------------------
type rx_sync_fsm_type is (
   LOST_SYNC_ST,  --! IDLE state of the FSM
   CHECK_SYNC_ST, --! Checking data to validate synchronization state
   READY_ST       --! Synchronization ok state
   );
---------------------------------------------------------
----- Signal declaration -----
---------------------------------------------------------
signal current_state                : rx_sync_fsm_type;                                    --! Current state of the Lane Initialization FSM
signal comma_det_PLWA_r             : std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! COMMA_DET_PLWA registered signal
signal data_rx_to_lcwd_i            : std_logic_vector(C_DATA_WIDTH-1 downto 0);          --! 64-bit data sent to lane_ctrl_word_detect
signal valid_k_charac_to_lcwd_i     : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags to lane_ctrl_word_detect
signal data_rdy_to_lcwd_i           : std_logic;                                           --! Data valid flag to lane_ctrl_word_detect
signal err_word_cnt                 : unsigned(2 downto 0);                                --! RXERR control word counter
signal err_word_x5                  : std_logic;                                           --! Flag indicates that err_word_cnt reaches 5
signal valid_symb                   : std_logic;                                           --! Flag indicates that a valid symbol is received
signal disp_invalid_err             : std_logic;                                           --! Flag indicates that a disparity error or an invalid symbol is detected

begin
---------------------------------------------------------
-----                   Assignation                 -----
---------------------------------------------------------
DATA_RX_PLRSF        <= data_rx_to_lcwd_i;
VALID_K_CHARAC_PLRSF <= valid_k_charac_to_lcwd_i;
DATA_RDY_PLRSF       <= data_rdy_to_lcwd_i;
---------------------------------------------------------
-----               Process                         -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_rx_sync_fsm_transition
--! Receiver word synchronization FSM transition process
---------------------------------------------------------
  p_rx_sync_fsm_transition : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      current_state              <= LOST_SYNC_ST;
      comma_det_PLWA_r        <= (others => '0');
    elsif rising_edge(CLK) then
      comma_det_PLWA_r        <= COMMA_DET_PLWA;
      case current_state is
        when LOST_SYNC_ST   =>  if COMMA_DET_PLWA /= std_logic_vector(to_unsigned(0, COMMA_DET_PLWA'length)) then -- when a Comma sequence is detected
                                  current_state  <= CHECK_SYNC_ST;
                                else
                                  current_state  <= LOST_SYNC_ST;
                                end if;
        when CHECK_SYNC_ST  =>  if (LANE_RESET = '1' or LANE_RESET_DL = '1') or RX_WORD_IS_ALIGNED_PLWA = '0' or err_word_x5 = '1' then
                                  current_state  <= LOST_SYNC_ST;
                                elsif valid_symb = '1' then
                                  current_state  <= READY_ST;
                                else
                                  current_state  <= CHECK_SYNC_ST;
                                end if;
        when READY_ST       =>  if (LANE_RESET = '1' or LANE_RESET_DL = '1') or RX_WORD_IS_ALIGNED_PLWA = '0' then
                                  current_state  <= LOST_SYNC_ST;
                                elsif disp_invalid_err= '1' then
                                  current_state  <= CHECK_SYNC_ST;
                                else
                                  current_state  <= READY_ST;
                                end if;
        when others         => current_state  <= LOST_SYNC_ST;
      end case;
    end if;
  end process p_rx_sync_fsm_transition;
---------------------------------------------------------
-- Process: p_rx_sync_action_on_state
--! Receiver word synchronization FSM actions on state process
---------------------------------------------------------
  p_rx_sync_action_on_state : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      data_rx_to_lcwd_i          <= (others => '0');
      valid_k_charac_to_lcwd_i   <= (others => '0');
      data_rdy_to_lcwd_i         <= '0';
      err_word_cnt               <= (others => '0');
      err_word_x5                <= '0';
      valid_symb                 <= '0';
      disp_invalid_err           <= '0';
    elsif rising_edge(CLK) then
      if current_state = LOST_SYNC_ST then
        err_word_cnt               <= (others => '0');
        err_word_x5                <= '0';
        data_rx_to_lcwd_i          <= C_RXERR_WORD & C_RXERR_WORD;
        valid_k_charac_to_lcwd_i   <= x"11";
        data_rdy_to_lcwd_i         <= '1';
      elsif current_state = CHECK_SYNC_ST then
        disp_invalid_err           <= '0';
        data_rx_to_lcwd_i          <= DATA_RX_PLWA;
        valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_PLWA;
        data_rdy_to_lcwd_i         <= '1';
        -- Alignment valid and error flag de-asserted
        if err_word_x5 = '0' and RX_WORD_IS_ALIGNED_PLWA= '1' then
          ---------------------------------------------------------
          -- Invalid character or disparity error treatment --
          ---------------------------------------------------------
          -- Error in each word of the data bus
          if (INVALID_CHAR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0") and (INVALID_CHAR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0")then
            data_rx_to_lcwd_i          <= C_RXERR_WORD & C_RXERR_WORD;
            valid_k_charac_to_lcwd_i   <= x"11";
            if err_word_cnt >= C_SYMB_X5 then
              err_word_x5   <= '1';
            elsif err_word_cnt < C_SYMB_X5 then
              err_word_cnt  <= err_word_cnt + 2;
              err_word_x5   <= '0';
            end if;
          -- Error in the first word (only) of the data bus
          elsif INVALID_CHAR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" then
            data_rx_to_lcwd_i          <= DATA_RX_PLWA(C_DATA_WIDTH-1 downto C_DATA_WIDTH/2) & C_RXERR_WORD;
            valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) & x"1";
            valid_symb                 <= '1';
            err_word_cnt               <= (others => '0');
            err_word_x5                <= '0';
          -- Error in the second word (only) of the data bus
          elsif INVALID_CHAR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" then
            data_rx_to_lcwd_i          <= C_RXERR_WORD & DATA_RX_PLWA(C_DATA_WIDTH/2-1 downto 0);
            valid_k_charac_to_lcwd_i   <= x"1" & VALID_K_CHARAC_PLWA(C_K_CHAR_WIDTH/2-1 downto 0);
            err_word_cnt               <= to_unsigned(1,err_word_cnt'length);
            err_word_x5                <= '0';
          -- No error
          else
            valid_symb    <= '1';
            err_word_cnt  <= (others => '0');
            err_word_x5   <= '0';
          end if;
        else
            data_rx_to_lcwd_i          <= C_RXERR_WORD & C_RXERR_WORD;
            valid_k_charac_to_lcwd_i   <= x"11";
            valid_symb                 <= '0';
        end if;
      elsif current_state = READY_ST then
        err_word_cnt               <= (others => '0');
        valid_symb                 <= '0';
        data_rx_to_lcwd_i          <= DATA_RX_PLWA;
        valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_PLWA;
        data_rdy_to_lcwd_i         <= '1';
        if RX_WORD_IS_ALIGNED_PLWA= '1' then
          ---------------------------------------------------------
          -- Invalid character or disparity error treatment --
          ---------------------------------------------------------
          -- Error in each word of the data bus
          if (INVALID_CHAR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0") and (INVALID_CHAR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0")then
            data_rx_to_lcwd_i          <= C_RXERR_WORD & C_RXERR_WORD;
            valid_k_charac_to_lcwd_i   <= x"11";
            disp_invalid_err           <= '1';
          -- Error in the first word (only) of the data bus
          elsif INVALID_CHAR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH/2-1 downto 0) /= x"0" then
            data_rx_to_lcwd_i          <= DATA_RX_PLWA(C_DATA_WIDTH-1 downto C_DATA_WIDTH/2) & C_RXERR_WORD;
            valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) & x"1";
            disp_invalid_err           <= '0';
          -- Error in the second word (only) of the data bus
          elsif INVALID_CHAR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" or DISPARITY_ERR_PLWA(C_K_CHAR_WIDTH-1 downto C_K_CHAR_WIDTH/2) /= x"0" then
            data_rx_to_lcwd_i          <= C_RXERR_WORD & DATA_RX_PLWA(C_DATA_WIDTH/2-1 downto 0);
            valid_k_charac_to_lcwd_i   <= x"1" & VALID_K_CHARAC_PLWA(C_K_CHAR_WIDTH/2-1 downto 0);
            disp_invalid_err           <= '1';
          else
            -- No error
            disp_invalid_err           <= '0';
          end if;
        else
          data_rx_to_lcwd_i          <= C_RXERR_WORD & C_RXERR_WORD;
          valid_k_charac_to_lcwd_i   <= x"11";
        end if;
      end if;
    end if;
  end process p_rx_sync_action_on_state;
end architecture rtl;
