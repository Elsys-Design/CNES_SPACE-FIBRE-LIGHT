// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_FP_INMUX_DEFINES_VH
`else
`define B_DSP_FP_INMUX_DEFINES_VH

// Look-up table parameters
//

`define DSP_FP_INMUX_ADDR_N  10
`define DSP_FP_INMUX_ADDR_SZ 32
`define DSP_FP_INMUX_DATA_SZ 64

// Attribute addresses
//

`define DSP_FP_INMUX__AREG    32'h00000000
`define DSP_FP_INMUX__AREG_SZ 32

`define DSP_FP_INMUX__FPA_PREG    32'h00000001
`define DSP_FP_INMUX__FPA_PREG_SZ 32

`define DSP_FP_INMUX__FPBREG    32'h00000002
`define DSP_FP_INMUX__FPBREG_SZ 32

`define DSP_FP_INMUX__FPDREG    32'h00000003
`define DSP_FP_INMUX__FPDREG_SZ 32

`define DSP_FP_INMUX__INMODEREG    32'h00000004
`define DSP_FP_INMUX__INMODEREG_SZ 32

`define DSP_FP_INMUX__IS_FPINMODE_INVERTED    32'h00000005
`define DSP_FP_INMUX__IS_FPINMODE_INVERTED_SZ 1

`define DSP_FP_INMUX__IS_RSTFPINMODE_INVERTED    32'h00000006
`define DSP_FP_INMUX__IS_RSTFPINMODE_INVERTED_SZ 1

`define DSP_FP_INMUX__LEGACY    32'h00000007
`define DSP_FP_INMUX__LEGACY_SZ 40

`define DSP_FP_INMUX__RESET_MODE    32'h00000008
`define DSP_FP_INMUX__RESET_MODE_SZ 40

`define DSP_FP_INMUX__USE_MULT    32'h00000009
`define DSP_FP_INMUX__USE_MULT_SZ 64

`endif  // B_DSP_FP_INMUX_DEFINES_VH