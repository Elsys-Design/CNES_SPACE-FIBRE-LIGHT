// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_CMPHY_OCTAD_DEFINES_VH
`else
`define B_CMPHY_OCTAD_DEFINES_VH

// Look-up table parameters
//

`define CMPHY_OCTAD_ADDR_N  205
`define CMPHY_OCTAD_ADDR_SZ 32
`define CMPHY_OCTAD_DATA_SZ 160

// Attribute addresses
//

`define CMPHY_OCTAD__ACC_FAST_LOCK    32'h00000000
`define CMPHY_OCTAD__ACC_FAST_LOCK_SZ 56

`define CMPHY_OCTAD__APBCLK_FREQ    32'h00000001
`define CMPHY_OCTAD__APBCLK_FREQ_SZ 9

`define CMPHY_OCTAD__CAL_DQS_SRC    32'h00000002
`define CMPHY_OCTAD__CAL_DQS_SRC_SZ 64

`define CMPHY_OCTAD__CAL_REFCLK_EN    32'h00000003
`define CMPHY_OCTAD__CAL_REFCLK_EN_SZ 2

`define CMPHY_OCTAD__CAL_VT_OFST_C    32'h00000004
`define CMPHY_OCTAD__CAL_VT_OFST_C_SZ 10

`define CMPHY_OCTAD__CAL_VT_OFST_EN    32'h00000005
`define CMPHY_OCTAD__CAL_VT_OFST_EN_SZ 56

`define CMPHY_OCTAD__CAL_VT_OFST_M0    32'h00000006
`define CMPHY_OCTAD__CAL_VT_OFST_M0_SZ 10

`define CMPHY_OCTAD__CAL_VT_OFST_M1    32'h00000007
`define CMPHY_OCTAD__CAL_VT_OFST_M1_SZ 10

`define CMPHY_OCTAD__CAL_VT_SRC    32'h00000008
`define CMPHY_OCTAD__CAL_VT_SRC_SZ 48

`define CMPHY_OCTAD__CLB_CLK_DBL_DCC    32'h00000009
`define CMPHY_OCTAD__CLB_CLK_DBL_DCC_SZ 3

`define CMPHY_OCTAD__CLK_SRC    32'h0000000a
`define CMPHY_OCTAD__CLK_SRC_SZ 1

`define CMPHY_OCTAD__CLOCK_FREQ    32'h0000000b
`define CMPHY_OCTAD__CLOCK_FREQ_SZ 13

`define CMPHY_OCTAD__CN_EXT_DISABLE    32'h0000000c
`define CMPHY_OCTAD__CN_EXT_DISABLE_SZ 40

`define CMPHY_OCTAD__CN_LEGACY    32'h0000000d
`define CMPHY_OCTAD__CN_LEGACY_SZ 40

`define CMPHY_OCTAD__CONTINUOUS_DQS    32'h0000000e
`define CMPHY_OCTAD__CONTINUOUS_DQS_SZ 40

`define CMPHY_OCTAD__CPHY_RX_EN_0    32'h0000000f
`define CMPHY_OCTAD__CPHY_RX_EN_0_SZ 40

`define CMPHY_OCTAD__CPHY_RX_EN_1    32'h00000010
`define CMPHY_OCTAD__CPHY_RX_EN_1_SZ 40

`define CMPHY_OCTAD__CPHY_TX_EN_0    32'h00000011
`define CMPHY_OCTAD__CPHY_TX_EN_0_SZ 40

`define CMPHY_OCTAD__CPHY_TX_EN_1    32'h00000012
`define CMPHY_OCTAD__CPHY_TX_EN_1_SZ 40

`define CMPHY_OCTAD__CTLE_OFST_CAL_0    32'h00000013
`define CMPHY_OCTAD__CTLE_OFST_CAL_0_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_1    32'h00000014
`define CMPHY_OCTAD__CTLE_OFST_CAL_1_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_2    32'h00000015
`define CMPHY_OCTAD__CTLE_OFST_CAL_2_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_3    32'h00000016
`define CMPHY_OCTAD__CTLE_OFST_CAL_3_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_4    32'h00000017
`define CMPHY_OCTAD__CTLE_OFST_CAL_4_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_5    32'h00000018
`define CMPHY_OCTAD__CTLE_OFST_CAL_5_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_6    32'h00000019
`define CMPHY_OCTAD__CTLE_OFST_CAL_6_SZ 128

`define CMPHY_OCTAD__CTLE_OFST_CAL_7    32'h0000001a
`define CMPHY_OCTAD__CTLE_OFST_CAL_7_SZ 128

`define CMPHY_OCTAD__DCC_CAL_RANGE    32'h0000001b
`define CMPHY_OCTAD__DCC_CAL_RANGE_SZ 12

`define CMPHY_OCTAD__DCC_CAL_TIME_SEL    32'h0000001c
`define CMPHY_OCTAD__DCC_CAL_TIME_SEL_SZ 152

`define CMPHY_OCTAD__DCC_CONV_RANGE    32'h0000001d
`define CMPHY_OCTAD__DCC_CONV_RANGE_SZ 12

`define CMPHY_OCTAD__DCC_CONV_TIME_SEL    32'h0000001e
`define CMPHY_OCTAD__DCC_CONV_TIME_SEL_SZ 160

`define CMPHY_OCTAD__DCC_RO_DLY0    32'h0000001f
`define CMPHY_OCTAD__DCC_RO_DLY0_SZ 9

`define CMPHY_OCTAD__DCC_RO_DLY1    32'h00000020
`define CMPHY_OCTAD__DCC_RO_DLY1_SZ 9

`define CMPHY_OCTAD__DCC_RO_DLY2    32'h00000021
`define CMPHY_OCTAD__DCC_RO_DLY2_SZ 9

`define CMPHY_OCTAD__DMC_APB_SEL    32'h00000022
`define CMPHY_OCTAD__DMC_APB_SEL_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_0    32'h00000023
`define CMPHY_OCTAD__DMC_BIT_SEL_0_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_1    32'h00000024
`define CMPHY_OCTAD__DMC_BIT_SEL_1_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_2    32'h00000025
`define CMPHY_OCTAD__DMC_BIT_SEL_2_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_3    32'h00000026
`define CMPHY_OCTAD__DMC_BIT_SEL_3_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_4    32'h00000027
`define CMPHY_OCTAD__DMC_BIT_SEL_4_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_5    32'h00000028
`define CMPHY_OCTAD__DMC_BIT_SEL_5_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_6    32'h00000029
`define CMPHY_OCTAD__DMC_BIT_SEL_6_SZ 40

`define CMPHY_OCTAD__DMC_BIT_SEL_7    32'h0000002a
`define CMPHY_OCTAD__DMC_BIT_SEL_7_SZ 40

`define CMPHY_OCTAD__DMC_CTL_SEL    32'h0000002b
`define CMPHY_OCTAD__DMC_CTL_SEL_SZ 40

`define CMPHY_OCTAD__DPHY_RX_EN_0    32'h0000002c
`define CMPHY_OCTAD__DPHY_RX_EN_0_SZ 40

`define CMPHY_OCTAD__DPHY_RX_EN_1    32'h0000002d
`define CMPHY_OCTAD__DPHY_RX_EN_1_SZ 40

`define CMPHY_OCTAD__DPHY_RX_EN_2    32'h0000002e
`define CMPHY_OCTAD__DPHY_RX_EN_2_SZ 40

`define CMPHY_OCTAD__DPHY_RX_EN_3    32'h0000002f
`define CMPHY_OCTAD__DPHY_RX_EN_3_SZ 40

`define CMPHY_OCTAD__DPHY_TX_EN_0    32'h00000030
`define CMPHY_OCTAD__DPHY_TX_EN_0_SZ 40

`define CMPHY_OCTAD__DPHY_TX_EN_1    32'h00000031
`define CMPHY_OCTAD__DPHY_TX_EN_1_SZ 40

`define CMPHY_OCTAD__DPHY_TX_EN_2    32'h00000032
`define CMPHY_OCTAD__DPHY_TX_EN_2_SZ 40

`define CMPHY_OCTAD__DPHY_TX_EN_3    32'h00000033
`define CMPHY_OCTAD__DPHY_TX_EN_3_SZ 40

`define CMPHY_OCTAD__DQS_MODE    32'h00000034
`define CMPHY_OCTAD__DQS_MODE_SZ 3

`define CMPHY_OCTAD__EN_CK90_CAL    32'h00000035
`define CMPHY_OCTAD__EN_CK90_CAL_SZ 40

`define CMPHY_OCTAD__EN_DCC_CAL    32'h00000036
`define CMPHY_OCTAD__EN_DCC_CAL_SZ 40

`define CMPHY_OCTAD__EN_FIX_DELAY_CAL    32'h00000037
`define CMPHY_OCTAD__EN_FIX_DELAY_CAL_SZ 40

`define CMPHY_OCTAD__EN_PRIMARY_DLL_CAL    32'h00000038
`define CMPHY_OCTAD__EN_PRIMARY_DLL_CAL_SZ 40

`define CMPHY_OCTAD__EN_SEQ_CAL    32'h00000039
`define CMPHY_OCTAD__EN_SEQ_CAL_SZ 40

`define CMPHY_OCTAD__FD_NORD    32'h0000003a
`define CMPHY_OCTAD__FD_NORD_SZ 1

`define CMPHY_OCTAD__GT_VT_SRC    32'h0000003b
`define CMPHY_OCTAD__GT_VT_SRC_SZ 64

`define CMPHY_OCTAD__GT_VT_SRC_OCTAD    32'h0000003c
`define CMPHY_OCTAD__GT_VT_SRC_OCTAD_SZ 48

`define CMPHY_OCTAD__HISTO_DELTA_ADJ    32'h0000003d
`define CMPHY_OCTAD__HISTO_DELTA_ADJ_SZ 13

`define CMPHY_OCTAD__HISTO_F0_TH    32'h0000003e
`define CMPHY_OCTAD__HISTO_F0_TH_SZ 10

`define CMPHY_OCTAD__HISTO_F1_TH    32'h0000003f
`define CMPHY_OCTAD__HISTO_F1_TH_SZ 10

`define CMPHY_OCTAD__HISTO_NO_RU    32'h00000040
`define CMPHY_OCTAD__HISTO_NO_RU_SZ 40

`define CMPHY_OCTAD__HISTO_NPI_NS    32'h00000041
`define CMPHY_OCTAD__HISTO_NPI_NS_SZ 7

`define CMPHY_OCTAD__HISTO_R0_TH    32'h00000042
`define CMPHY_OCTAD__HISTO_R0_TH_SZ 10

`define CMPHY_OCTAD__HISTO_R1_TH    32'h00000043
`define CMPHY_OCTAD__HISTO_R1_TH_SZ 10

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_0    32'h00000044
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_0_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_1    32'h00000045
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_1_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_2    32'h00000046
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_2_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_3    32'h00000047
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_3_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_4    32'h00000048
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_4_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_5    32'h00000049
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_5_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_6    32'h0000004a
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_6_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_7    32'h0000004b
`define CMPHY_OCTAD__IBUF_DIS_EXT_SRC_7_SZ 40

`define CMPHY_OCTAD__IBUF_DIS_SRC_0    32'h0000004c
`define CMPHY_OCTAD__IBUF_DIS_SRC_0_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_1    32'h0000004d
`define CMPHY_OCTAD__IBUF_DIS_SRC_1_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_2    32'h0000004e
`define CMPHY_OCTAD__IBUF_DIS_SRC_2_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_3    32'h0000004f
`define CMPHY_OCTAD__IBUF_DIS_SRC_3_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_4    32'h00000050
`define CMPHY_OCTAD__IBUF_DIS_SRC_4_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_5    32'h00000051
`define CMPHY_OCTAD__IBUF_DIS_SRC_5_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_6    32'h00000052
`define CMPHY_OCTAD__IBUF_DIS_SRC_6_SZ 64

`define CMPHY_OCTAD__IBUF_DIS_SRC_7    32'h00000053
`define CMPHY_OCTAD__IBUF_DIS_SRC_7_SZ 64

`define CMPHY_OCTAD__LEG_F_HISTO_E    32'h00000054
`define CMPHY_OCTAD__LEG_F_HISTO_E_SZ 40

`define CMPHY_OCTAD__LEG_F_LGY_E    32'h00000055
`define CMPHY_OCTAD__LEG_F_LGY_E_SZ 40

`define CMPHY_OCTAD__MIPI_ALPRX_EN_M    32'h00000056
`define CMPHY_OCTAD__MIPI_ALPRX_EN_M_SZ 40

`define CMPHY_OCTAD__MIPI_ALPRX_EN_S    32'h00000057
`define CMPHY_OCTAD__MIPI_ALPRX_EN_S_SZ 40

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_0    32'h00000058
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_0_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_1    32'h00000059
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_1_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_2    32'h0000005a
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_2_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_3    32'h0000005b
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_3_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_4    32'h0000005c
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_4_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_5    32'h0000005d
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_5_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_6    32'h0000005e
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_6_SZ 10

`define CMPHY_OCTAD__NQTR_DELAY_VALUE_7    32'h0000005f
`define CMPHY_OCTAD__NQTR_DELAY_VALUE_7_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_0    32'h00000060
`define CMPHY_OCTAD__O_DELAY_VALUE_0_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_1    32'h00000061
`define CMPHY_OCTAD__O_DELAY_VALUE_1_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_2    32'h00000062
`define CMPHY_OCTAD__O_DELAY_VALUE_2_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_3    32'h00000063
`define CMPHY_OCTAD__O_DELAY_VALUE_3_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_4    32'h00000064
`define CMPHY_OCTAD__O_DELAY_VALUE_4_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_5    32'h00000065
`define CMPHY_OCTAD__O_DELAY_VALUE_5_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_6    32'h00000066
`define CMPHY_OCTAD__O_DELAY_VALUE_6_SZ 10

`define CMPHY_OCTAD__O_DELAY_VALUE_7    32'h00000067
`define CMPHY_OCTAD__O_DELAY_VALUE_7_SZ 10

`define CMPHY_OCTAD__PDL_CASCADE    32'h00000068
`define CMPHY_OCTAD__PDL_CASCADE_SZ 40

`define CMPHY_OCTAD__PDL_HISTOGRAM_MODE    32'h00000069
`define CMPHY_OCTAD__PDL_HISTOGRAM_MODE_SZ 56

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_0    32'h0000006a
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_0_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_1    32'h0000006b
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_1_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_2    32'h0000006c
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_2_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_3    32'h0000006d
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_3_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_4    32'h0000006e
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_4_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_5    32'h0000006f
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_5_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_6    32'h00000070
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_6_SZ 10

`define CMPHY_OCTAD__PQTR_DELAY_VALUE_7    32'h00000071
`define CMPHY_OCTAD__PQTR_DELAY_VALUE_7_SZ 10

`define CMPHY_OCTAD__PRIMARY_DLL_CONFIG    32'h00000072
`define CMPHY_OCTAD__PRIMARY_DLL_CONFIG_SZ 48

`define CMPHY_OCTAD__RIUCLK_DBLR_BYPASS    32'h00000073
`define CMPHY_OCTAD__RIUCLK_DBLR_BYPASS_SZ 40

`define CMPHY_OCTAD__RIU_CLK_DBL_DCC    32'h00000074
`define CMPHY_OCTAD__RIU_CLK_DBL_DCC_SZ 3

`define CMPHY_OCTAD__ROUTETHRU_0    32'h00000075
`define CMPHY_OCTAD__ROUTETHRU_0_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_1    32'h00000076
`define CMPHY_OCTAD__ROUTETHRU_1_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_2    32'h00000077
`define CMPHY_OCTAD__ROUTETHRU_2_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_3    32'h00000078
`define CMPHY_OCTAD__ROUTETHRU_3_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_4    32'h00000079
`define CMPHY_OCTAD__ROUTETHRU_4_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_5    32'h0000007a
`define CMPHY_OCTAD__ROUTETHRU_5_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_6    32'h0000007b
`define CMPHY_OCTAD__ROUTETHRU_6_SZ 40

`define CMPHY_OCTAD__ROUTETHRU_7    32'h0000007c
`define CMPHY_OCTAD__ROUTETHRU_7_SZ 40

`define CMPHY_OCTAD__RXFIFO_MODE_0    32'h0000007d
`define CMPHY_OCTAD__RXFIFO_MODE_0_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_1    32'h0000007e
`define CMPHY_OCTAD__RXFIFO_MODE_1_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_2    32'h0000007f
`define CMPHY_OCTAD__RXFIFO_MODE_2_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_3    32'h00000080
`define CMPHY_OCTAD__RXFIFO_MODE_3_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_4    32'h00000081
`define CMPHY_OCTAD__RXFIFO_MODE_4_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_5    32'h00000082
`define CMPHY_OCTAD__RXFIFO_MODE_5_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_6    32'h00000083
`define CMPHY_OCTAD__RXFIFO_MODE_6_SZ 48

`define CMPHY_OCTAD__RXFIFO_MODE_7    32'h00000084
`define CMPHY_OCTAD__RXFIFO_MODE_7_SZ 48

`define CMPHY_OCTAD__RXFIFO_WRCLK_SEL    32'h00000085
`define CMPHY_OCTAD__RXFIFO_WRCLK_SEL_SZ 32

`define CMPHY_OCTAD__RXOFST_CAL_START    32'h00000086
`define CMPHY_OCTAD__RXOFST_CAL_START_SZ 4

`define CMPHY_OCTAD__RXOFST_END_CODE    32'h00000087
`define CMPHY_OCTAD__RXOFST_END_CODE_SZ 8

`define CMPHY_OCTAD__RXOFST_EN_BIN_SRCH    32'h00000088
`define CMPHY_OCTAD__RXOFST_EN_BIN_SRCH_SZ 1

`define CMPHY_OCTAD__RXOFST_EN_HIST_SRCH    32'h00000089
`define CMPHY_OCTAD__RXOFST_EN_HIST_SRCH_SZ 1

`define CMPHY_OCTAD__RXOFST_EN_LIN_SRCH    32'h0000008a
`define CMPHY_OCTAD__RXOFST_EN_LIN_SRCH_SZ 1

`define CMPHY_OCTAD__RXOFST_EXTEND_OFSC_RANGE    32'h0000008b
`define CMPHY_OCTAD__RXOFST_EXTEND_OFSC_RANGE_SZ 40

`define CMPHY_OCTAD__RXOFST_EXTRANGE_STEPSIZE    32'h0000008c
`define CMPHY_OCTAD__RXOFST_EXTRANGE_STEPSIZE_SZ 7

`define CMPHY_OCTAD__RXOFST_LIN_SRCH_RANGE    32'h0000008d
`define CMPHY_OCTAD__RXOFST_LIN_SRCH_RANGE_SZ 5

`define CMPHY_OCTAD__RXOFST_LIN_SRCH_STEPSIZE    32'h0000008e
`define CMPHY_OCTAD__RXOFST_LIN_SRCH_STEPSIZE_SZ 2

`define CMPHY_OCTAD__RXOFST_NUM_SAMPLES    32'h0000008f
`define CMPHY_OCTAD__RXOFST_NUM_SAMPLES_SZ 11

`define CMPHY_OCTAD__RXOFST_SETTELE_INTERVAL    32'h00000090
`define CMPHY_OCTAD__RXOFST_SETTELE_INTERVAL_SZ 5

`define CMPHY_OCTAD__RXOFST_START_CODE    32'h00000091
`define CMPHY_OCTAD__RXOFST_START_CODE_SZ 8

`define CMPHY_OCTAD__RXOFST_THRESHOLD    32'h00000092
`define CMPHY_OCTAD__RXOFST_THRESHOLD_SZ 8

`define CMPHY_OCTAD__RX_CLOCK_ALIGN    32'h00000093
`define CMPHY_OCTAD__RX_CLOCK_ALIGN_SZ 152

`define CMPHY_OCTAD__RX_DATA_WIDTH    32'h00000094
`define CMPHY_OCTAD__RX_DATA_WIDTH_SZ 5

`define CMPHY_OCTAD__RX_PATH_RESET    32'h00000095
`define CMPHY_OCTAD__RX_PATH_RESET_SZ 56

`define CMPHY_OCTAD__SA_OFST_CAL_0    32'h00000096
`define CMPHY_OCTAD__SA_OFST_CAL_0_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_1    32'h00000097
`define CMPHY_OCTAD__SA_OFST_CAL_1_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_2    32'h00000098
`define CMPHY_OCTAD__SA_OFST_CAL_2_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_3    32'h00000099
`define CMPHY_OCTAD__SA_OFST_CAL_3_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_4    32'h0000009a
`define CMPHY_OCTAD__SA_OFST_CAL_4_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_5    32'h0000009b
`define CMPHY_OCTAD__SA_OFST_CAL_5_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_6    32'h0000009c
`define CMPHY_OCTAD__SA_OFST_CAL_6_SZ 112

`define CMPHY_OCTAD__SA_OFST_CAL_7    32'h0000009d
`define CMPHY_OCTAD__SA_OFST_CAL_7_SZ 112

`define CMPHY_OCTAD__SEQ_DIS_0    32'h0000009e
`define CMPHY_OCTAD__SEQ_DIS_0_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_1    32'h0000009f
`define CMPHY_OCTAD__SEQ_DIS_1_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_2    32'h000000a0
`define CMPHY_OCTAD__SEQ_DIS_2_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_3    32'h000000a1
`define CMPHY_OCTAD__SEQ_DIS_3_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_4    32'h000000a2
`define CMPHY_OCTAD__SEQ_DIS_4_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_5    32'h000000a3
`define CMPHY_OCTAD__SEQ_DIS_5_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_6    32'h000000a4
`define CMPHY_OCTAD__SEQ_DIS_6_SZ 40

`define CMPHY_OCTAD__SEQ_DIS_7    32'h000000a5
`define CMPHY_OCTAD__SEQ_DIS_7_SZ 40

`define CMPHY_OCTAD__SEQ_DONE_MASK    32'h000000a6
`define CMPHY_OCTAD__SEQ_DONE_MASK_SZ 4

`define CMPHY_OCTAD__SEQ_DQS_CENTER    32'h000000a7
`define CMPHY_OCTAD__SEQ_DQS_CENTER_SZ 2

`define CMPHY_OCTAD__SEQ_HISTROGRAM_MODE    32'h000000a8
`define CMPHY_OCTAD__SEQ_HISTROGRAM_MODE_SZ 56

`define CMPHY_OCTAD__SIM_VERSION    32'h000000a9
`define CMPHY_OCTAD__SIM_VERSION_SZ 2

`define CMPHY_OCTAD__SLEW_MODE    32'h000000aa
`define CMPHY_OCTAD__SLEW_MODE_SZ 40

`define CMPHY_OCTAD__TBYTE_CTL_0    32'h000000ab
`define CMPHY_OCTAD__TBYTE_CTL_0_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_1    32'h000000ac
`define CMPHY_OCTAD__TBYTE_CTL_1_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_2    32'h000000ad
`define CMPHY_OCTAD__TBYTE_CTL_2_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_3    32'h000000ae
`define CMPHY_OCTAD__TBYTE_CTL_3_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_4    32'h000000af
`define CMPHY_OCTAD__TBYTE_CTL_4_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_5    32'h000000b0
`define CMPHY_OCTAD__TBYTE_CTL_5_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_6    32'h000000b1
`define CMPHY_OCTAD__TBYTE_CTL_6_SZ 64

`define CMPHY_OCTAD__TBYTE_CTL_7    32'h000000b2
`define CMPHY_OCTAD__TBYTE_CTL_7_SZ 64

`define CMPHY_OCTAD__TX_DATA_WIDTH    32'h000000b3
`define CMPHY_OCTAD__TX_DATA_WIDTH_SZ 5

`define CMPHY_OCTAD__TX_FIFO_PD_OFFSET    32'h000000b4
`define CMPHY_OCTAD__TX_FIFO_PD_OFFSET_SZ 3

`define CMPHY_OCTAD__TX_FIFO_SYNC_BYPASS    32'h000000b5
`define CMPHY_OCTAD__TX_FIFO_SYNC_BYPASS_SZ 40

`define CMPHY_OCTAD__TX_INIT_0    32'h000000b6
`define CMPHY_OCTAD__TX_INIT_0_SZ 40

`define CMPHY_OCTAD__TX_INIT_1    32'h000000b7
`define CMPHY_OCTAD__TX_INIT_1_SZ 40

`define CMPHY_OCTAD__TX_INIT_2    32'h000000b8
`define CMPHY_OCTAD__TX_INIT_2_SZ 40

`define CMPHY_OCTAD__TX_INIT_3    32'h000000b9
`define CMPHY_OCTAD__TX_INIT_3_SZ 40

`define CMPHY_OCTAD__TX_INIT_4    32'h000000ba
`define CMPHY_OCTAD__TX_INIT_4_SZ 40

`define CMPHY_OCTAD__TX_INIT_5    32'h000000bb
`define CMPHY_OCTAD__TX_INIT_5_SZ 40

`define CMPHY_OCTAD__TX_INIT_6    32'h000000bc
`define CMPHY_OCTAD__TX_INIT_6_SZ 40

`define CMPHY_OCTAD__TX_INIT_7    32'h000000bd
`define CMPHY_OCTAD__TX_INIT_7_SZ 40

`define CMPHY_OCTAD__TX_INIT_T    32'h000000be
`define CMPHY_OCTAD__TX_INIT_T_SZ 40

`define CMPHY_OCTAD__VTC_NOT_SPD    32'h000000bf
`define CMPHY_OCTAD__VTC_NOT_SPD_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_0    32'h000000c0
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_0_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_1    32'h000000c1
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_1_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_2    32'h000000c2
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_2_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_3    32'h000000c3
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_3_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_4    32'h000000c4
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_4_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_5    32'h000000c5
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_5_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_6    32'h000000c6
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_6_SZ 40

`define CMPHY_OCTAD__WREN_CS_OVERRIDE_7    32'h000000c7
`define CMPHY_OCTAD__WREN_CS_OVERRIDE_7_SZ 40

`define CMPHY_OCTAD__WR_CTL_MUXSEL    32'h000000c8
`define CMPHY_OCTAD__WR_CTL_MUXSEL_SZ 8

`define CMPHY_OCTAD__WR_DQ0_MUXSEL    32'h000000c9
`define CMPHY_OCTAD__WR_DQ0_MUXSEL_SZ 8

`define CMPHY_OCTAD__WR_DQ1_MUXSEL    32'h000000ca
`define CMPHY_OCTAD__WR_DQ1_MUXSEL_SZ 8

`define CMPHY_OCTAD__WR_EN0_MUXSEL    32'h000000cb
`define CMPHY_OCTAD__WR_EN0_MUXSEL_SZ 8

`define CMPHY_OCTAD__WR_EN1_MUXSEL    32'h000000cc
`define CMPHY_OCTAD__WR_EN1_MUXSEL_SZ 8

`endif  // B_CMPHY_OCTAD_DEFINES_VH