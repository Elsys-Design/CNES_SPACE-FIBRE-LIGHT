library IEEE;
use IEEE.std_logic_1164.all;

library phy_plus_lane_lib;
 use phy_plus_lane_lib.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

library interlayer_lib;
use interlayer_lib.all;

entity spacefibre_light_top_ip is
   port (
          RST_N                            : in  std_logic;                            --! global reset
      CLK                              : in  std_logic;                            --! Main clock
      CLK_TX                           : out  std_logic;                           --! Clock generated by manufacturer IP
      RST_TXCLK_N                      : out  std_logic;                           --! Reset clock generated by manufacturer IP
      -- CLK GTY signals
      CLK_GTY                          : in std_logic;                             --! GTY dedicated clock
      -- FROM/TO Outside
      TX_POS                           : out std_logic;                            --! Positive LVDS serial data send
      TX_NEG                           : out std_logic;                            --! Negative LVDS serial data send
      RX_POS                           : in  std_logic;                            --! Positive LVDS serial data received
      RX_NEG                           : in  std_logic;                            --! Negative LVDS serial data received
      ----------------------- Data-Link layer signals -----------------------


      -- virtual channels spacefibre axistream
      AXIS_ACLK_RX_DL        :  in  std_logic_vector(8 downto 0);
      AXIS_ACLK_TX_DL        :  in  std_logic_vector(8 downto 0);
      AXIS_ARSTN_RX_DL       :  in  std_logic_vector(8 downto 0);
      AXIS_ARSTN_TX_DL       :  in  std_logic_vector(8 downto 0);
      AXIS_TDATA_TX_DL_0     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_1     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_2     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_3     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_4     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_5     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_6     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_7     :  in  std_logic_vector(31 downto 0);
      AXIS_TDATA_TX_DL_8     :  in  std_logic_vector(31 downto 0);
      AXIS_TLAST_TX_DL       :  in  std_logic_vector(8 downto 0);
      AXIS_TREADY_RX_DL      :  in  std_logic_vector(8 downto 0);
      AXIS_TUSER_TX_DL_0     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_1     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_2     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_3     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_4     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_5     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_6     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_7     :  in  std_logic_vector(3 downto 0);
      AXIS_TUSER_TX_DL_8     :  in  std_logic_vector(3 downto 0);
      AXIS_TVALID_TX_DL      :  in  std_logic_vector(8 downto 0);

      AXIS_TDATA_RX_DL_0    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_1    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_2    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_3    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_4    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_5    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_6    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_7    :  out  std_logic_vector(31 downto 0);
      AXIS_TDATA_RX_DL_8    :  out  std_logic_vector(31 downto 0);
      AXIS_TLAST_RX_DL       :  out  std_logic_vector(8 downto 0);
      AXIS_TREADY_TX_DL      :  out  std_logic_vector(8 downto 0);
      AXIS_TUSER_RX_DL_0    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_1    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_2    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_3    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_4    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_5    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_6    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_7    :  out  std_logic_vector(3 downto 0);
      AXIS_TUSER_RX_DL_8    :  out  std_logic_vector(3 downto 0);
      AXIS_TVALID_RX_DL      :  out  std_logic_vector(8 downto 0);

      CURRENT_TIME_SLOT_NW             : in  std_logic_vector(7 downto 0);         --! Current time slot

   -- Parameters signals
      INTERFACE_RESET                  : in  std_logic;                            --! Reset the link and all configuration register of the Data Link layer
      LINK_RESET                       : in  std_logic;                            --! Reset the link
      NACK_RST_EN                      : in  std_logic;                            --! Enable automatic link reset on NACK reception
      NACK_RST_MODE                    : in  std_logic;                            --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
      PAUSE_VC                         : in  std_logic_vector(8 downto 0);         --! Pause the corresponding virtual channel after the end of current transmission
      CONTINUOUS_VC                    : in  std_logic_vector(7 downto 0);         --! Enable the corresponding virtual channel continuous mode
      -- Status signals
      SEQ_NUMBER_TX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in transmission
      SEQ_NUMBER_RX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in reception
      CREDIT_VC                        : out std_logic_vector(7 downto 0);          --! Indicates if each corresponding far-end input buffer has credit
      INPUT_BUF_OVF_VC                 : out std_logic_vector(7 downto 0); --! Indicates input buffer overflow
      FCT_CREDIT_OVERFLOW              : out std_logic_vector(7 downto 0);          --! Indicates overflow of each corresponding input buffer
      CRC_LONG_ERROR                   : out std_logic;                             --! CRC long error
      CRC_SHORT_ERROR                  : out std_logic;                             --! CRC short error
      FRAME_ERROR                      : out std_logic;                             --! Frame error
      SEQUENCE_ERROR                   : out std_logic;                             --! Sequence error
      FAR_END_LINK_RESET               : out std_logic;                             --! Far-end link reset status
      FRAME_FINISHED                   : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel finished emitting a frame
      FRAME_TX                         : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel is emitting a frame
      DATA_COUNTER_TX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data transmitted in last frame emitted
      DATA_COUNTER_RX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data received in last frame received
      ACK_COUNTER_TX                   : out std_logic_vector(2 downto 0);          --! ACK counter TX
      NACK_COUNTER_TX                  : out std_logic_vector(2 downto 0);          --! NACK counter TX
      FCT_COUNTER_TX                   : out std_logic_vector(3 downto 0);          --! FCT counter TX
      ACK_COUNTER_RX                   : out std_logic_vector(2 downto 0);          --! ACK counter RX
      NACK_COUNTER_RX                  : out std_logic_vector(2 downto 0);          --! NACK counter RX
      FCT_COUNTER_RX                   : out std_logic_vector(3 downto 0);          --! FCT counter RX
      FULL_COUNTER_RX                  : out std_logic_vector(1 downto 0);          --! FULL counter RX
      RETRY_COUNTER_RX                 : out std_logic_vector(1 downto 0);          --! RETRY counter RX
      CURRENT_TIME_SLOT                : out std_logic_vector(7 downto 0);          --! Current time slot
      RESET_PARAM                      : out std_logic;                             --! Reset parameters register command
      LINK_RST_ASSERTED                : out std_logic;                             --! Link reset status
      NACK_SEQ_NUM                     : out std_logic_vector(7 downto 0);          --! NACK Seq_num received
      ACK_SEQ_NUM                      : out std_logic_vector(7 downto 0);          --! ACK Seq_num received
      DATA_PULSE_RX                    : out std_logic;                             --! Data received pulse signal
      ACK_PULSE_RX                     : out std_logic;                             --! ACK received pulse signal
      NACK_PULSE_RX                    : out std_logic;                             --! NACK received pulse signal
      FCT_PULSE_RX                     : out std_logic;                             --! FCT received pulse signal
      FULL_PULSE_RX                    : out std_logic;                             --! FULL received pulse signal
      RETRY_PULSE_RX                   : out std_logic;                             --! RETRY received pulse signal
      ----------------------- Phy + Lane layer signals -----------------------
      -- -- Interface injector
      ENABLE_INJ                       : in std_logic;                              --! Enable injector command
      DATA_TX_INJ                      : in  std_logic_vector(31 downto 00);        --! Data parallel to be send from injector
      CAPABILITY_TX_INJ                : in  std_logic_vector(07 downto 00);        --! Capability send on TX link in INIT3 control word from injector
      NEW_DATA_TX_INJ                  : in  std_logic;                             --! Flag to write data in FIFO TX from injetor
      VALID_K_CHARAC_TX_INJ            : in  std_logic_vector(03 downto 00);        --! K charachter valid in the 32-bit DATA_TX_INJ vector
      FIFO_TX_FULL_INJ                 : out   std_logic;                           --! Flag full of the FIFO TX to the injector
      LANE_RESET_INJ                   : in  std_logic;                             --! Lane Reset command from Injector
      -- -- Interface spy
      ENABLE_SPY                       : in std_logic;                              --! Enable Spy read command
      FIFO_RX_RD_EN_SPY                : in  std_logic;                             --! FiFo RX read enable flag from the spy
      DATA_RX_SPY                      : out std_logic_vector(31 downto 00);        --! 32-bit Data parallel to be received to the spy
      FIFO_RX_EMPTY_SPY                : out std_logic;                             --! FiFo RX empty flag to the spy
      FIFO_RX_DATA_VALID_SPY           : out std_logic;                             --! FiFo RX data valid flag to the spy
      VALID_K_CHARAC_RX_SPY            : out std_logic_vector(03 downto 00);        --! 4-bit valid K character flags to the spy
      -- Paramter and Status signals
      LANE_START                       : in  std_logic;                             --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                             --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                             --! Asserts or de-asserts LaneReset for the lane
      PARALLEL_LOOPBACK_EN             : in  std_logic;                             --! Enables or disables the parallel loopback for the lane
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);        --! In case of error, pauses communication
      NEAR_END_SERIAL_LB_EN            : in  std_logic;                             --! Enables or disables the near-end serial loopback for the lane
      FAR_END_SERIAL_LB_EN             : in  std_logic;                             --! Enables or disables the far-end serial loopback for the lane
      LANE_STATE                       : out std_logic_vector(03 downto 00);        --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);        --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic;                             --! Overflow flag of the RX_ERROR_CNT
      LOSS_SIGNAL                      : out std_logic;                             --! Set when no signal is received on RX link
      FAR_END_CAPA                     : out std_logic_vector(07 downto 00);        --! RX Capabilities field (INT3 flags)
      RX_POLARITY                      : out std_logic                              --! Set when the receiver polarity is inverted
   );
end entity spacefibre_light_top_ip;

architecture rtl of spacefibre_light_top_ip is
 constant G_VC_NUM                         : integer := 8 ;
 
        -- Component declaration for spacefibre_light_top
        component spacefibre_light_top is
            generic(
                G_VC_NUM                         : integer := 8                                    --! Number of virtual channel
                );
             port (
  RST_N                            : in  std_logic;                            --! global reset
      CLK                              : in  std_logic;                            --! Main clock
      CLK_TX                           : out  std_logic;                           --! Clock generated by manufacturer IP
      RST_TXCLK_N                      : out  std_logic;                           --! Reset clock generated by manufacturer IP
      -- CLK GTY signals
      CLK_GTY                          : in std_logic;                             --! GTY dedicated clock
      -- FROM/TO Outside
      TX_POS                           : out std_logic;                            --! Positive LVDS serial data send
      TX_NEG                           : out std_logic;                            --! Negative LVDS serial data send
      RX_POS                           : in  std_logic;                            --! Positive LVDS serial data received
      RX_NEG                           : in  std_logic;                            --! Negative LVDS serial data received
      ----------------------- Data-Link layer signals -----------------------
      -- Discret signals
      AXIS_ARSTN_TX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Active-low asynchronous reset signals for each virtual channel (VC) in the TX path
      AXIS_ACLK_TX_DL                  : in  std_logic_vector(G_VC_NUM downto 0);  --! Clock signals for each VC in the TX path
      AXIS_TREADY_TX_DL                : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates that the data link layer is ready to accept data on each VC
      AXIS_TDATA_TX_DL                 : in  vc_data_array(G_VC_NUM downto 0);     --! Data signals from the network layer to the data link layer for each VC
      AXIS_TUSER_TX_DL                 : in  vc_k_array(G_VC_NUM downto 0);        --! Sideband information (e.g., control or metadata) from the network layer to the data link layer for each VC
      AXIS_TLAST_TX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates the last transfer in a packet/transaction on each VC
      AXIS_TVALID_TX_DL                : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates that valid data is available on the TX data bus for each VC
      AXIS_ARSTN_RX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Active-low asynchronous reset signals for each VC in the RX path
      AXIS_ACLK_RX_DL                  : in  std_logic_vector(G_VC_NUM downto 0);  --! Clock signals for each VC in the RX path
      AXIS_TREADY_RX_DL                : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates that the network layer is ready to receive data on each VC
      AXIS_TDATA_RX_DL                 : out vc_data_array(G_VC_NUM downto 0);     --! Data signals from the data link layer to the network layer for each VC
      AXIS_TUSER_RX_DL                 : out vc_k_array(G_VC_NUM downto 0);        --! Sideband information from the data link layer to the network layer for each VC
      AXIS_TLAST_RX_DL                 : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates the last transfer in a packet/transaction on each VC
      AXIS_TVALID_RX_DL                : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates that valid data is available on the RX data bus for each VC
      CURRENT_TIME_SLOT_NW             : in  std_logic_vector(7 downto 0);         --! Current time slot
      -- Paramters signals
      INTERFACE_RESET                  : in  std_logic;                            --! Reset the link and all configuration register of the Data Link layer
      LINK_RESET                       : in  std_logic;                            --! Reset the link
      NACK_RST_EN                      : in  std_logic;                            --! Enable automatic link reset on NACK reception
      NACK_RST_MODE                    : in  std_logic;                            --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
      PAUSE_VC                         : in  std_logic_vector(8 downto 0);         --! Pause the corresponding virtual channel after the end of current transmission
      CONTINUOUS_VC                    : in  std_logic_vector(7 downto 0);         --! Enable the corresponding virtual channel continuous mode
      -- Status signals
      SEQ_NUMBER_TX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in transmission
      SEQ_NUMBER_RX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in reception
      CREDIT_VC                        : out std_logic_vector(7 downto 0);          --! Indicates if each corresponding far-end input buffer has credit
      INPUT_BUF_OVF_VC                 : out std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates input buffer overflow
      FCT_CREDIT_OVERFLOW              : out std_logic_vector(7 downto 0);          --! Indicates overflow of each corresponding input buffer
      CRC_LONG_ERROR                   : out std_logic;                             --! CRC long error
      CRC_SHORT_ERROR                  : out std_logic;                             --! CRC short error
      FRAME_ERROR                      : out std_logic;                             --! Frame error
      SEQUENCE_ERROR                   : out std_logic;                             --! Sequence error
      FAR_END_LINK_RESET               : out std_logic;                             --! Far-end link reset status
      FRAME_FINISHED                   : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel finished emitting a frame
      FRAME_TX                         : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel is emitting a frame
      DATA_COUNTER_TX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data transmitted in last frame emitted
      DATA_COUNTER_RX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data received in last frame received
      ACK_COUNTER_TX                   : out std_logic_vector(2 downto 0);          --! ACK counter TX
      NACK_COUNTER_TX                  : out std_logic_vector(2 downto 0);          --! NACK counter TX
      FCT_COUNTER_TX                   : out std_logic_vector(3 downto 0);          --! FCT counter TX
      ACK_COUNTER_RX                   : out std_logic_vector(2 downto 0);          --! ACK counter RX
      NACK_COUNTER_RX                  : out std_logic_vector(2 downto 0);          --! NACK counter RX
      FCT_COUNTER_RX                   : out std_logic_vector(3 downto 0);          --! FCT counter RX
      FULL_COUNTER_RX                  : out std_logic_vector(1 downto 0);          --! FULL counter RX
      RETRY_COUNTER_RX                 : out std_logic_vector(1 downto 0);          --! RETRY counter RX
      CURRENT_TIME_SLOT                : out std_logic_vector(7 downto 0);          --! Current time slot
      RESET_PARAM                      : out std_logic;                             --! Reset parameters register command
      LINK_RST_ASSERTED                : out std_logic;                             --! Link reset status
      NACK_SEQ_NUM                     : out std_logic_vector(7 downto 0);          --! NACK Seq_num received
      ACK_SEQ_NUM                      : out std_logic_vector(7 downto 0);          --! ACK Seq_num received
      DATA_PULSE_RX                    : out std_logic;                             --! Data received pulse signal
      ACK_PULSE_RX                     : out std_logic;                             --! ACK received pulse signal
      NACK_PULSE_RX                    : out std_logic;                             --! NACK received pulse signal
      FCT_PULSE_RX                     : out std_logic;                             --! FCT received pulse signal
      FULL_PULSE_RX                    : out std_logic;                             --! FULL received pulse signal
      RETRY_PULSE_RX                   : out std_logic;                             --! RETRY received pulse signal
      ----------------------- Phy + Lane layer signals -----------------------
      -- -- Interface injector
      ENABLE_INJ                       : in std_logic;                              --! Enable injector command
      DATA_TX_INJ                      : in  std_logic_vector(31 downto 00);        --! Data parallel to be send from injector
      CAPABILITY_TX_INJ                : in  std_logic_vector(07 downto 00);        --! Capability send on TX link in INIT3 control word from injector
      NEW_DATA_TX_INJ                  : in  std_logic;                             --! Flag to write data in FIFO TX from injetor
      VALID_K_CHARAC_TX_INJ            : in  std_logic_vector(03 downto 00);        --! K charachter valid in the 32-bit DATA_TX_INJ vector
      FIFO_TX_FULL_INJ                 : out   std_logic;                           --! Flag full of the FIFO TX to the injector
      LANE_RESET_INJ                   : in  std_logic;                             --! Lane Reset command from Injector
      -- -- Interface spy
      ENABLE_SPY                       : in std_logic;                              --! Enable Spy read command
      FIFO_RX_RD_EN_SPY                : in  std_logic;                             --! FiFo RX read enable flag from the spy
      DATA_RX_SPY                      : out std_logic_vector(31 downto 00);        --! 32-bit Data parallel to be received to the spy
      FIFO_RX_EMPTY_SPY                : out std_logic;                             --! FiFo RX empty flag to the spy
      FIFO_RX_DATA_VALID_SPY           : out std_logic;                             --! FiFo RX data valid flag to the spy
      VALID_K_CHARAC_RX_SPY            : out std_logic_vector(03 downto 00);        --! 4-bit valid K character flags to the spy
      -- Paramter and Status signals
      LANE_START                       : in  std_logic;                             --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                             --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                             --! Asserts or de-asserts LaneReset for the lane
      PARALLEL_LOOPBACK_EN             : in  std_logic;                             --! Enables or disables the parallel loopback for the lane
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);        --! In case of error, pauses communication
      NEAR_END_SERIAL_LB_EN            : in  std_logic;                             --! Enables or disables the near-end serial loopback for the lane
      FAR_END_SERIAL_LB_EN             : in  std_logic;                             --! Enables or disables the far-end serial loopback for the lane
      LANE_STATE                       : out std_logic_vector(03 downto 00);        --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);        --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic;                             --! Overflow flag of the RX_ERROR_CNT
      LOSS_SIGNAL                      : out std_logic;                             --! Set when no signal is received on RX link
      FAR_END_CAPA                     : out std_logic_vector(07 downto 00);        --! RX Capabilities field (INT3 flags)
      RX_POLARITY                      : out std_logic                              --! Set when the receiver polarity is inverted
   );
        end component;
        

begin
spacefibre_light_top_inst: spacefibre_light_top
   generic map (G_VC_NUM=>G_VC_NUM)
   port map (
      -- Input Ports - Single Bit
      AUTOSTART                         => AUTOSTART,                       
      CLK                               => CLK,                             
      CLK_GTY                           => CLK_GTY,                         
      ENABLE_INJ                        => ENABLE_INJ,                      
      ENABLE_SPY                        => ENABLE_SPY,                      
      FAR_END_SERIAL_LB_EN              => FAR_END_SERIAL_LB_EN,            
      FIFO_RX_RD_EN_SPY                 => FIFO_RX_RD_EN_SPY,               
      INTERFACE_RESET                   => INTERFACE_RESET,                 
      LANE_RESET                        => LANE_RESET,                      
      LANE_RESET_INJ                    => LANE_RESET_INJ,                  
      LANE_START                        => LANE_START,                      
      LINK_RESET                        => LINK_RESET,                      
      NACK_RST_EN                       => NACK_RST_EN,                     
      NACK_RST_MODE                     => NACK_RST_MODE,                   
      NEAR_END_SERIAL_LB_EN             => NEAR_END_SERIAL_LB_EN,           
      NEW_DATA_TX_INJ                   => NEW_DATA_TX_INJ,                 
      PARALLEL_LOOPBACK_EN              => PARALLEL_LOOPBACK_EN,            
      RST_N                             => RST_N,                           
      RX_NEG                            => RX_NEG,                          
      RX_POS                            => RX_POS,                          
      -- Input Ports - Busses
      AXIS_ACLK_RX_DL(8 downto 0)       => AXIS_ACLK_RX_DL(8 downto 0),     
      AXIS_ACLK_TX_DL(8 downto 0)       => AXIS_ACLK_TX_DL(8 downto 0),     
      AXIS_ARSTN_RX_DL(8 downto 0)      => AXIS_ARSTN_RX_DL(8 downto 0),    
      AXIS_ARSTN_TX_DL(8 downto 0)      => AXIS_ARSTN_TX_DL(8 downto 0),    
      AXIS_TDATA_TX_DL(0)(31 downto 0)  => AXIS_TDATA_TX_DL_0(31 downto 0),
      AXIS_TDATA_TX_DL(1)(31 downto 0)  => AXIS_TDATA_TX_DL_1(31 downto 0),
      AXIS_TDATA_TX_DL(2)(31 downto 0)  => AXIS_TDATA_TX_DL_2(31 downto 0),
      AXIS_TDATA_TX_DL(3)(31 downto 0)  => AXIS_TDATA_TX_DL_3(31 downto 0),
      AXIS_TDATA_TX_DL(4)(31 downto 0)  => AXIS_TDATA_TX_DL_4(31 downto 0),
      AXIS_TDATA_TX_DL(5)(31 downto 0)  => AXIS_TDATA_TX_DL_5(31 downto 0),
      AXIS_TDATA_TX_DL(6)(31 downto 0)  => AXIS_TDATA_TX_DL_6(31 downto 0),
      AXIS_TDATA_TX_DL(7)(31 downto 0)  => AXIS_TDATA_TX_DL_7(31 downto 0),
      AXIS_TDATA_TX_DL(8)(31 downto 0)  => AXIS_TDATA_TX_DL_8(31 downto 0),
      AXIS_TLAST_TX_DL(8 downto 0)      => AXIS_TLAST_TX_DL(8 downto 0),    
      AXIS_TREADY_RX_DL(8 downto 0)     => AXIS_TREADY_RX_DL(8 downto 0),   
      AXIS_TUSER_TX_DL(0)(3 downto 0)   => AXIS_TUSER_TX_DL_0(3 downto 0), 
      AXIS_TUSER_TX_DL(1)(3 downto 0)   => AXIS_TUSER_TX_DL_1(3 downto 0), 
      AXIS_TUSER_TX_DL(2)(3 downto 0)   => AXIS_TUSER_TX_DL_2(3 downto 0), 
      AXIS_TUSER_TX_DL(3)(3 downto 0)   => AXIS_TUSER_TX_DL_3(3 downto 0), 
      AXIS_TUSER_TX_DL(4)(3 downto 0)   => AXIS_TUSER_TX_DL_4(3 downto 0), 
      AXIS_TUSER_TX_DL(5)(3 downto 0)   => AXIS_TUSER_TX_DL_5(3 downto 0), 
      AXIS_TUSER_TX_DL(6)(3 downto 0)   => AXIS_TUSER_TX_DL_6(3 downto 0), 
      AXIS_TUSER_TX_DL(7)(3 downto 0)   => AXIS_TUSER_TX_DL_7(3 downto 0), 
      AXIS_TUSER_TX_DL(8)(3 downto 0)   => AXIS_TUSER_TX_DL_8(3 downto 0), 
      AXIS_TVALID_TX_DL(8 downto 0)     => AXIS_TVALID_TX_DL(8 downto 0),   
      CAPABILITY_TX_INJ(7 downto 0)     => CAPABILITY_TX_INJ(7 downto 0),   
      CONTINUOUS_VC(7 downto 0)         => CONTINUOUS_VC(7 downto 0),       
      CURRENT_TIME_SLOT_NW(7 downto 0)  => CURRENT_TIME_SLOT_NW(7 downto 0),
      DATA_TX_INJ(31 downto 0)          => DATA_TX_INJ(31 downto 0),        
      PAUSE_VC(8 downto 0)              => PAUSE_VC(8 downto 0),            
      STANDBY_REASON(7 downto 0)        => STANDBY_REASON(7 downto 0),      
      VALID_K_CHARAC_TX_INJ(3 downto 0) => VALID_K_CHARAC_TX_INJ(3 downto 0),
      -- Output Ports - Single Bit
      ACK_PULSE_RX                      => ACK_PULSE_RX,                    
      CLK_TX                            => CLK_TX,                          
      CRC_LONG_ERROR                    => CRC_LONG_ERROR,                  
      CRC_SHORT_ERROR                   => CRC_SHORT_ERROR,                 
      DATA_PULSE_RX                     => DATA_PULSE_RX,                   
      FAR_END_LINK_RESET                => FAR_END_LINK_RESET,              
      FCT_PULSE_RX                      => FCT_PULSE_RX,                    
      FIFO_RX_DATA_VALID_SPY            => FIFO_RX_DATA_VALID_SPY,          
      FIFO_RX_EMPTY_SPY                 => FIFO_RX_EMPTY_SPY,               
      FIFO_TX_FULL_INJ                  => FIFO_TX_FULL_INJ,                
      FRAME_ERROR                       => FRAME_ERROR,                     
      FULL_PULSE_RX                     => FULL_PULSE_RX,                   
      LINK_RST_ASSERTED                 => LINK_RST_ASSERTED,               
      LOSS_SIGNAL                       => LOSS_SIGNAL,                     
      NACK_PULSE_RX                     => NACK_PULSE_RX,                   
      RESET_PARAM                       => RESET_PARAM,                     
      RETRY_PULSE_RX                    => RETRY_PULSE_RX,                  
      RST_TXCLK_N                       => RST_TXCLK_N,                     
      RX_ERROR_OVF                      => RX_ERROR_OVF,                    
      RX_POLARITY                       => RX_POLARITY,                     
      SEQUENCE_ERROR                    => SEQUENCE_ERROR,                  
      TX_NEG                            => TX_NEG,                          
      TX_POS                            => TX_POS,                          
      -- Output Ports - Busses
      ACK_COUNTER_RX(2 downto 0)        => ACK_COUNTER_RX(2 downto 0),      
      ACK_COUNTER_TX(2 downto 0)        => ACK_COUNTER_TX(2 downto 0),      
      ACK_SEQ_NUM(7 downto 0)           => ACK_SEQ_NUM(7 downto 0),         
      AXIS_TDATA_RX_DL(0)(31 downto 0)  => AXIS_TDATA_RX_DL_0(31 downto 0),
      AXIS_TDATA_RX_DL(1)(31 downto 0)  => AXIS_TDATA_RX_DL_1(31 downto 0),
      AXIS_TDATA_RX_DL(2)(31 downto 0)  => AXIS_TDATA_RX_DL_2(31 downto 0),
      AXIS_TDATA_RX_DL(3)(31 downto 0)  => AXIS_TDATA_RX_DL_3(31 downto 0),
      AXIS_TDATA_RX_DL(4)(31 downto 0)  => AXIS_TDATA_RX_DL_4(31 downto 0),
      AXIS_TDATA_RX_DL(5)(31 downto 0)  => AXIS_TDATA_RX_DL_5(31 downto 0),
      AXIS_TDATA_RX_DL(6)(31 downto 0)  => AXIS_TDATA_RX_DL_6(31 downto 0),
      AXIS_TDATA_RX_DL(7)(31 downto 0)  => AXIS_TDATA_RX_DL_7(31 downto 0),
      AXIS_TDATA_RX_DL(8)(31 downto 0)  => AXIS_TDATA_RX_DL_8(31 downto 0),
      AXIS_TLAST_RX_DL(8 downto 0)      => AXIS_TLAST_RX_DL(8 downto 0),    
      AXIS_TREADY_TX_DL(8 downto 0)     => AXIS_TREADY_TX_DL(8 downto 0),   
      AXIS_TUSER_RX_DL(0)(3 downto 0)   => AXIS_TUSER_RX_DL_0(3 downto 0), 
      AXIS_TUSER_RX_DL(1)(3 downto 0)   => AXIS_TUSER_RX_DL_1(3 downto 0), 
      AXIS_TUSER_RX_DL(2)(3 downto 0)   => AXIS_TUSER_RX_DL_2(3 downto 0), 
      AXIS_TUSER_RX_DL(3)(3 downto 0)   => AXIS_TUSER_RX_DL_3(3 downto 0), 
      AXIS_TUSER_RX_DL(4)(3 downto 0)   => AXIS_TUSER_RX_DL_4(3 downto 0), 
      AXIS_TUSER_RX_DL(5)(3 downto 0)   => AXIS_TUSER_RX_DL_5(3 downto 0), 
      AXIS_TUSER_RX_DL(6)(3 downto 0)   => AXIS_TUSER_RX_DL_6(3 downto 0), 
      AXIS_TUSER_RX_DL(7)(3 downto 0)   => AXIS_TUSER_RX_DL_7(3 downto 0), 
      AXIS_TUSER_RX_DL(8)(3 downto 0)   => AXIS_TUSER_RX_DL_8(3 downto 0), 
      AXIS_TVALID_RX_DL(8 downto 0)     => AXIS_TVALID_RX_DL(8 downto 0),   
      CREDIT_VC(7 downto 0)             => CREDIT_VC(7 downto 0),           
      CURRENT_TIME_SLOT(7 downto 0)     => CURRENT_TIME_SLOT(7 downto 0),   
      DATA_COUNTER_RX(6 downto 0)       => DATA_COUNTER_RX(6 downto 0),     
      DATA_COUNTER_TX(6 downto 0)       => DATA_COUNTER_TX(6 downto 0),     
      DATA_RX_SPY(31 downto 0)          => DATA_RX_SPY(31 downto 0),        
      FAR_END_CAPA(7 downto 0)          => FAR_END_CAPA(7 downto 0),        
      FCT_COUNTER_RX(3 downto 0)        => FCT_COUNTER_RX(3 downto 0),      
      FCT_COUNTER_TX(3 downto 0)        => FCT_COUNTER_TX(3 downto 0),      
      FCT_CREDIT_OVERFLOW(7 downto 0)   => FCT_CREDIT_OVERFLOW(7 downto 0), 
      FRAME_FINISHED(8 downto 0)        => FRAME_FINISHED(8 downto 0),      
      FRAME_TX(8 downto 0)              => FRAME_TX(8 downto 0),            
      FULL_COUNTER_RX(1 downto 0)       => FULL_COUNTER_RX(1 downto 0),     
      INPUT_BUF_OVF_VC(7 downto 0)      => INPUT_BUF_OVF_VC(7 downto 0),    
      LANE_STATE(3 downto 0)            => LANE_STATE(3 downto 0),          
      NACK_COUNTER_RX(2 downto 0)       => NACK_COUNTER_RX(2 downto 0),     
      NACK_COUNTER_TX(2 downto 0)       => NACK_COUNTER_TX(2 downto 0),     
      NACK_SEQ_NUM(7 downto 0)          => NACK_SEQ_NUM(7 downto 0),        
      RETRY_COUNTER_RX(1 downto 0)      => RETRY_COUNTER_RX(1 downto 0),    
      RX_ERROR_CNT(7 downto 0)          => RX_ERROR_CNT(7 downto 0),        
      SEQ_NUMBER_RX(7 downto 0)         => SEQ_NUMBER_RX(7 downto 0),       
      SEQ_NUMBER_TX(7 downto 0)         => SEQ_NUMBER_TX(7 downto 0),       
      VALID_K_CHARAC_RX_SPY(3 downto 0) => VALID_K_CHARAC_RX_SPY(3 downto 0)
      -- InOut Ports - Single Bit
      -- InOut Ports - Busses
   );
end architecture rtl;