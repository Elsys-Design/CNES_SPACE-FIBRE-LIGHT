// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_ODELAYE3_DEFINES_VH
`else
`define B_ODELAYE3_DEFINES_VH

// Look-up table parameters
//

`define ODELAYE3_ADDR_N  10
`define ODELAYE3_ADDR_SZ 32
`define ODELAYE3_DATA_SZ 152

// Attribute addresses
//

`define ODELAYE3__CASCADE    32'h00000000
`define ODELAYE3__CASCADE_SZ 96

`define ODELAYE3__DELAY_FORMAT    32'h00000001
`define ODELAYE3__DELAY_FORMAT_SZ 40

`define ODELAYE3__DELAY_TYPE    32'h00000002
`define ODELAYE3__DELAY_TYPE_SZ 64

`define ODELAYE3__DELAY_VALUE    32'h00000003
`define ODELAYE3__DELAY_VALUE_SZ 32

`define ODELAYE3__IS_CLK_INVERTED    32'h00000004
`define ODELAYE3__IS_CLK_INVERTED_SZ 1

`define ODELAYE3__IS_RST_INVERTED    32'h00000005
`define ODELAYE3__IS_RST_INVERTED_SZ 1

`define ODELAYE3__REFCLK_FREQUENCY    32'h00000006
`define ODELAYE3__REFCLK_FREQUENCY_SZ 64

`define ODELAYE3__SIM_DEVICE    32'h00000007
`define ODELAYE3__SIM_DEVICE_SZ 152

`define ODELAYE3__SIM_VERSION    32'h00000008
`define ODELAYE3__SIM_VERSION_SZ 64

`define ODELAYE3__UPDATE_MODE    32'h00000009
`define ODELAYE3__UPDATE_MODE_SZ 48

`endif  // B_ODELAYE3_DEFINES_VH