----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description : This module describe the Lane_init_FSM function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
use phy_plus_lane_lib.all;

entity lane_init_fsm is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP
      -- FROM/TO Data-link layer
      LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer.

      -- RX signals
      NO_SIGNAL                        : in  std_logic;                       --! Flag no signal are received
      RX_NEW_WORD                      : in  std_logic;                       --! Flag new word has been received
      DETECTED_INIT1                   : in  std_logic;                       --! Flag INIT1 control word rxed
      DETECTED_INIT2                   : in  std_logic;                       --! Flag INIT2 control word rxed
      DETECTED_INIT3                   : in  std_logic;                       --! Flag INIT3 control word rxed
      DETECTED_INV_INIT1               : in  std_logic;                       --! Flag INV_INIT1 control word rxed
      DETECTED_INV_INIT2               : in  std_logic;                       --! Flag INV_INIT2 control word rxed
      DETECTED_RXERR_WORD              : in  std_logic;                       --! Flag RXERR detected
      DETECTED_LOSS_SIGNAL             : in  std_logic;                       --! Flag LOSS_SINGAL control word detected
      DETECTED_STANDBY                 : in  std_logic;                       --! Flag STANDBY control word detected
      COMMA_K287_RXED                  : in  std_logic;                       --! Flag Comma K28.7 has been received
      RECEIVER_DISABLED                : out std_logic;                       --! flag to enabled RX function of HSSL IP
      CDR                              : out std_logic;                       --! Flag to enabled CDR function of HSSL IP
      SEND_RXERR                       : out std_logic;                       --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
      INVERT_RX_BITS                   : out std_logic;                       --! Flag to Invert rx bit received
      NO_SIGNAL_DETECTION_ENABLED      : out std_logic;                       --! Flag to enable the no signal function

      -- TX signals
      STANDBY_SIGNAL_X32               : in  std_logic;                       --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32                  : in  std_logic;                       --! Flag LOST_SIGNAL control word has been send x32
      TRANSMITTER_DISABLED             : out std_logic;                       --! flag to enabled TX fonction of HSSL IP
      SEND_INIT1_CTRL_WORD             : out std_logic;                       --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD             : out std_logic;                       --! Flag to send control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD             : out std_logic;                       --! Flag to send control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA               : out std_logic;                       --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS       : out std_logic;                       --! Flag to send STANDBY control word x32
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   : out std_logic;                       --! Flag to send LOSS_SIGNAL control word x32
      LOST_CAUSE                       : out std_logic_vector(01 downto 00);  --! Flag to indicate the reason of the LOST_SIGNAL

      -- PARAMETERS and STATUS
      LANE_START                       : in  std_logic;                       --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                       --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                       --! Asserts or de-asserts LaneReset for the lane
      LANE_STATE                       : out std_logic_vector(03 downto 00);  --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic                        --! Overflow flag of the RX_ERROR_CNT
   );
end lane_init_fsm;

architecture rtl of lane_init_fsm is

----------------------------- Declaration signals -----------------------------

-- Lane Initialisation FSM transition conditions process
   -- Type
type lane_init_fsm_type is (
   CLEAR_LINE_ST,                                                                --! Reset state
   DISABLED_ST,                                                                  --! Disabled TX and RX State
   WAIT_ST,                                                                      --! Waiting State
   STARTED_ST,                                                                   --! Configuration INIT1 State
   INVERT_RX_POLARITY_ST,                                                        --! Invert RX polarity in case of detection invert control words
   CONNECTING_ST,                                                                --! Configuration INIT2 State
   CONNECTED_ST,                                                                 --! Configuration INIT3 State
   ACTIVE_ST,                                                                    --! Transmission Data State
   LOSS_OF_SIGNAL_ST,                                                            --! Error state loss of signal
   PREPARE_STANDBY_ST                                                            --! Error state standby
   );
   -- Signals
signal current_state                : lane_init_fsm_type;                        --! Current state of the Lane Initialisation FSM
signal current_state_r              : lane_init_fsm_type;                        --! Current state registered

-- Lane Initialisation FSM action on state process -------------------------------------------------------------
   -- Constants
constant C_2US_AT_150MHZ            : unsigned(08 downto 00) := "1" & x"2B";     --! 300 x 6.667ns = 2us
   -- Signals
signal clear_line_cnt               : unsigned(08 downto 00);                    --! 2us counter
signal clear_line_done              : std_logic;                                 --! Flag indicates that clear_line_cnt reaches C_2US_AT_150MHZ
signal cdr_i                        : std_logic;                                 --! CDR enable command
signal enable_init_cnt              : std_logic;                                 --! enable timeout initialisation counter flag

--RX words counter process -------------------------------------------------------------------------------------
   -- Constants
constant C_MAX_RX_WORDS             : unsigned(13 downto 00) := "11" & x"FFF";   --! 16384 words received
   -- Signals
signal rx_words_cnt                 : unsigned(13 downto 00);                    --! Number of words received counter
signal rx_new_word_r                : std_logic;                                 --! RX_NEW_WORD registered signal

-- RX error counter process ------------------------------------------------------------------------------------
   -- Constants
constant C_MAX_RXERR_CTRL_WORDS     : unsigned(07 downto 00) := x"FF";           --! 256 RXERR control words received
   -- Signals
signal rx_error_cnt_i               : unsigned(07 downto 00);                    --! RXERR control words counter
signal rx_error_cnt_ovf_i           : std_logic;                                 --! RXERR overflow flag
signal detected_rxerr_word_r        : std_logic;                                 --! DETECTED_RXERR_WORD registered signal

-- init_timeout_counter process --------------------------------------------------------------------------------
   -- Constants
constant C_32US_AT_150MHZ           : unsigned(12 downto 00) := "1" & x"2C0";    --! 4497 x 6.667ns = 32us
   -- Signals
signal init_timeout_cnt             : unsigned(12 downto 00);                    --! Initialisation timeout counter
signal init_timeout_reaches         : std_logic;                                 --! Flag indicates that init_timeout_cnt reaches C_32US_AT_150MHZ

-- Detection 3 consecutive LOST_SIGNAL process -----------------------------------------------------------------
   -- Signals
signal loss_signal_x3_cnt           : unsigned(01 downto 00);                    --! Detection of consecutive LOSS_SIGNAL control words received
signal lost_signal_x3               : std_logic;                                 --! Flag indicates that 3 consecutive LOSS_SIGNAL control word has been received

-- Detection 3 consecutive STANDBY process ---------------------------------------------------------------------
   -- Signals
signal standby_signal_x3_cnt        : unsigned(01 downto 00);                    --! Detection of consecutive STANDBY control words received
signal standby_signal_x3            : std_logic;                                 --! Flag indicates that 3 consecutive STANDBY control word has been received

-- INIT1 detection process -------------------------------------------------------------------------------------
   -- Signals
signal inv_init1_rxed_cnt           : unsigned(01 downto 00);                    --! Detection of the inversed INIT1 counter
signal init1_rxed                   : std_logic;                                 --! Flag indicates that an INIT1 control word has been received
signal init1_rxed_r                 : std_logic;                                 --! init1_rxed registered signal
signal inv_init1_rxed_x3            : std_logic;                                 --! Flag indicates that inv_init1_rxed_cnt reaches 3
signal detected_init1_r             : std_logic;                                 --! DETECTED_INIT1 registered signal
signal detected_inv_init1_r         : std_logic;                                 --! DETECTED_INV_INIT1 registered signal

-- INIT2 detection process ------------------------------------------------------------------------------------
   -- Signals
signal init2_rxed_cnt               : unsigned(01 downto 00);                    --! Detection of the INIT1 counter
signal inv_init2_rxed_cnt           : unsigned(01 downto 00);                    --! Detection of the inversed INIT1 counter
signal init2_rxed_x3                : std_logic;                                 --! Flag indicates that x3 INIT2 control word has been received
signal inv_init2_rxed_x3            : std_logic;                                 --! Flag indicates that inv_init2_rxed_cnt reaches 3
signal init2_rxed                   : std_logic;                                 --! Flag indicates that INIT2 control word has been received
signal detected_init2_r             : std_logic;                                 --! DETECTED_INIT2 registered signal
signal detected_inv_init2_r         : std_logic;                                 --! DETECTED_INV_INIT2 registered signal

-- INIT3 detection process ------------------------------------------------------------------------------------
   -- Signals
signal init3_rxed_cnt               : unsigned(01 downto 00);                    --! Detection of the INIT3 counter
signal init3_rxed_x3                : std_logic;                                 --! Flag indicates that x3 INIT3 control word has been received
signal detected_init3_r             : std_logic;                                 --! DETECTED_INIT3 registered signal
signal comma_k287_rxed_r            : std_logic;                                 --! COMMA_K287_RXED registered signal

-- Process for detection the reception of 1023 words including the reception of at least on INIT1 or INIT2 without RXERR control words
   -- Constants
constant C_1023_WORDS               : unsigned(09 downto 00) := "11" & x"FF";    --! 1023 words received in STARTED_ST or INVERT_RX_POLARITY_ST
   -- Signals
signal rxed_1023_word_cnt           : unsigned(09 downto 00);                    --! Counter of received words
signal rxed_1023_word               : std_logic;                                 --! Flag indicates that rxed_1023_word_cnt reaches C_1023_WORDS



begin

-------------------------------------------------------------------------------------------
   -- Lane Initialisation FSM transition conditions process
   p_fsm_lane_init_transition : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         current_state     <= CLEAR_LINE_ST;
         current_state_r   <= CLEAR_LINE_ST;

      elsif rising_edge(CLK) then

         current_state_r   <= current_state;

         case current_state is

            when CLEAR_LINE_ST         => if clear_line_done = '1' then          -- when 2u counter reaches
                                             current_state  <= DISABLED_ST;
                                          else
                                             current_state  <= CLEAR_LINE_ST;
                                          end if;

            when DISABLED_ST           => if LANE_RESET = '1' or LANE_RESET_DL = '1' then -- When a soft reset appears
                                             current_state  <= CLEAR_LINE_ST;
                                          elsif LANE_START = '1' or AUTOSTART = '1' then  -- When a start command is detected
                                             current_state  <= WAIT_ST;
                                          else
                                             current_state  <= DISABLED_ST;
                                          end if;

            when WAIT_ST               => if LANE_RESET = '1' or LANE_RESET_DL = '1' then -- When a soft reset appears
                                             current_state  <= CLEAR_LINE_ST;
                                          elsif LANE_START = '0' and AUTOSTART = '0' then -- When a start command is not detected
                                             current_state  <= DISABLED_ST;
                                          elsif LANE_START = '1' or NO_SIGNAL = '0' then  -- When a start command is detected or signal is received
                                             current_state  <= STARTED_ST;
                                          else
                                             current_state  <= WAIT_ST;
                                          end if;

            when STARTED_ST            => if (lost_signal_x3 = '1' or standby_signal_x3 = '1') or init_timeout_reaches = '1' or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state <= CLEAR_LINE_ST;
                                          elsif inv_init1_rxed_x3 = '1' or inv_init2_rxed_x3 = '1' then
                                             current_state  <= INVERT_RX_POLARITY_ST;
                                          elsif rxed_1023_word = '1' then
                                             current_state  <= CONNECTING_ST;
                                          else
                                             current_state  <= STARTED_ST;
                                          end if;

            when INVERT_RX_POLARITY_ST => if NO_SIGNAL = '1' or init_timeout_reaches = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state  <= CLEAR_LINE_ST;
                                          elsif rxed_1023_word = '1' then
                                             current_state  <= CONNECTING_ST;
                                          else
                                             current_state  <= INVERT_RX_POLARITY_ST;
                                          end if;

            when CONNECTING_ST         => if NO_SIGNAL = '1' or init_timeout_reaches = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state  <= CLEAR_LINE_ST;
                                          elsif init2_rxed_x3 = '1' or init3_rxed_x3 = '1' then
                                             current_state  <= CONNECTED_ST;
                                          else
                                             current_state  <= CONNECTING_ST;
                                          end if;

            when CONNECTED_ST          => if NO_SIGNAL = '1' or init_timeout_reaches = '1' or comma_k287_rxed_r = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state  <= CLEAR_LINE_ST;
                                          elsif init3_rxed_x3 = '1' then
                                             current_state  <= ACTIVE_ST;
                                          else
                                             current_state  <= CONNECTED_ST;
                                          end if;

            when ACTIVE_ST             => if (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state <= CLEAR_LINE_ST;
                                          elsif LANE_START = '0' and AUTOSTART = '0' then
                                             current_state  <= PREPARE_STANDBY_ST;
                                          elsif init1_rxed = '1' or NO_SIGNAL = '1' or rx_error_cnt_ovf_i = '1' then
                                             current_state  <= LOSS_OF_SIGNAL_ST;
                                          else
                                             current_state  <= ACTIVE_ST;
                                          end if;

            when LOSS_OF_SIGNAL_ST     => if LOST_SIGNAL_X32 = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state <= CLEAR_LINE_ST;
                                          else
                                             current_state  <= LOSS_OF_SIGNAL_ST;
                                          end if;

            when PREPARE_STANDBY_ST    => if STANDBY_SIGNAL_X32 = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET = '1' or LANE_RESET_DL = '1' then
                                             current_state <= CLEAR_LINE_ST;
                                          else
                                             current_state  <= PREPARE_STANDBY_ST;
                                          end if;

            when others                => current_state  <= CLEAR_LINE_ST;

         end case;
      end if;
   end process p_fsm_lane_init_transition;

-------------------------------------------------------------------------------------------
   -- Lane Initialisation FSM action on state process
   p_comb_state : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         clear_line_cnt                      <= (others => '0');  -- Counter 2us of CLEAR_LINE_ST
         clear_line_done                     <= '0';              -- End condition of CLEAR_LINE_ST
         RECEIVER_DISABLED                   <= '1';              -- Receiver Disable
         TRANSMITTER_DISABLED                <= '1';              -- Transmitter Disabled
         cdr_i                               <= '0';              -- CDR Disabled
         SEND_INIT1_CTRL_WORD                <= '0';              -- stop send INIT1 control word following by 64 pseudo-random data words
         SEND_INIT2_CTRL_WORD                <= '0';              -- stop INIT2 control word following by 64 pseudo-random data words
         SEND_INIT3_CTRL_WORD                <= '0';              -- stop INIT3 control word following by 64 pseudo-random data words
         enable_init_cnt                     <= '0';              -- enable timeout initialisation counter
         INVERT_RX_BITS                      <= '0';              -- do not invert received bits
         ENABLE_TRANSM_DATA                  <= '0';              -- enable transimission data and control word from data-link layer
         SEND_32_STANDBY_CTRL_WORDS          <= '0';              -- stop 32 STANDBY control words
         SEND_32_LOSS_SIGNAL_CTRL_WORDS      <= '0';              -- stop 32 LOSS_SIGNAL control words
         NO_SIGNAL_DETECTION_ENABLED         <= '0';              -- No_signal detection function disabled
         LANE_STATE                          <= (others => '0');  -- Status of the Lane Init FSM
         LOST_CAUSE                          <= (others => '0');  -- LOST_SIGNAL reason

      elsif rising_edge(CLK) then

         if current_state = CLEAR_LINE_ST then

            LANE_STATE                       <= x"0"; -- Status of the FSM
            RECEIVER_DISABLED                <= '1';  -- Receiver Disable
            TRANSMITTER_DISABLED             <= '1';  -- Transmitter Disabled
            cdr_i                            <= '0';  -- CDR Disabled
            SEND_INIT1_CTRL_WORD             <= '0';  -- Send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '0';  -- Send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '0';  -- Send INIT3 control word following by 64 pseudo-random data words
            enable_init_cnt                  <= '0';  -- disable timeout initialisation counter
            INVERT_RX_BITS                   <= '0';  -- do not invert received bits
            ENABLE_TRANSM_DATA               <= '0';  -- disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS       <= '0';  -- Send 32 STANDBY control words
            SEND_32_LOSS_SIGNAL_CTRL_WORDS   <= '0';  -- Send 32 LOSS_SIGNAL control words
            NO_SIGNAL_DETECTION_ENABLED      <= '0';  -- No_signal detection function disabled
            LOST_CAUSE                       <= "00"; -- Reset

            -- Start counter 2us
            if clear_line_cnt >= C_2US_AT_150MHZ then
               clear_line_done   <= '1';              -- End condition of CLEAR_LINE_ST
            else
               clear_line_cnt    <= clear_line_cnt+1; -- Increment to 1 2us counter
               clear_line_done   <= '0';              -- Reset flag
            end if;

         elsif current_state = DISABLED_ST then

            clear_line_cnt                   <= (others => '0');  -- Reset 2us counter to 0
            LANE_STATE                       <= x"1"; -- Status of the FSM
            clear_line_done                  <= '0';  -- Reset 2us flag
            TRANSMITTER_DISABLED             <= '1';  -- Transmitter Disabled
            RECEIVER_DISABLED                <= '1';  -- Receiver Disabled
            cdr_i                            <= '0';  -- CDR Disabled

         elsif current_state = WAIT_ST then

            LANE_STATE                       <= x"2";
            RECEIVER_DISABLED                <= '0';  -- Receiver Enabled
            TRANSMITTER_DISABLED             <= '1';  -- Transmitter Disabled
            cdr_i                            <= '0';  -- CDR Disabled
            NO_SIGNAL_DETECTION_ENABLED      <= '1';  -- No_signal detection function enabled

         elsif current_state = STARTED_ST then

            LANE_STATE                       <= x"3"; -- Status of the FSM
            enable_init_cnt                  <= '1';  -- enable timeout initialisation counter
            TRANSMITTER_DISABLED             <= '0';  -- Transmitter Enable
            cdr_i                            <= '1';  -- CDR Enable
            SEND_INIT1_CTRL_WORD             <= '1';  -- send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = INVERT_RX_POLARITY_ST then

            LANE_STATE                       <= x"4"; -- Status of the FSM
            TRANSMITTER_DISABLED             <= '0';  -- Transmitter Enable
            cdr_i                            <= '1';  -- CDR Enable
            INVERT_RX_BITS                   <= '1';  -- invert received bits
            SEND_INIT1_CTRL_WORD             <= '1';  -- send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = CONNECTING_ST then

            LANE_STATE                       <= x"5";
            SEND_INIT1_CTRL_WORD             <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '1';  -- send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = CONNECTED_ST then

            LANE_STATE                       <= x"6"; -- Status of the FSM
            SEND_INIT1_CTRL_WORD             <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '1';  -- send INIT3 control word following by 64 pseudo-random data words

         elsif current_state = ACTIVE_ST then

            LANE_STATE                       <= x"7"; -- Status of the FSM
            SEND_INIT1_CTRL_WORD             <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD             <= '0';  -- send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD             <= '0';  -- send INIT3 control word following by 64 pseudo-random data words
            enable_init_cnt                  <= '0';  -- disable timeout initialisation counter
            ENABLE_TRANSM_DATA               <= '1';  -- enable transimission data and control word from data-link layer

         elsif current_state = PREPARE_STANDBY_ST then

            LANE_STATE                       <= x"8"; -- Status of the FSM
            ENABLE_TRANSM_DATA               <= '0';  -- Disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS       <= '1';  -- send 32 STANDBY control words

         elsif current_state = LOSS_OF_SIGNAL_ST then

            LANE_STATE                       <= x"9"; -- Status of the FSM
            ENABLE_TRANSM_DATA               <= '0';  -- Disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS       <= '0';  -- stop 32 STANDBY control words
            SEND_32_LOSS_SIGNAL_CTRL_WORDS   <= '1';  -- send 32 LOSS_SIGNAL control words

            -- Reason of the LOST_SIGNAL
            if init1_rxed_r = '1' then
               LOST_CAUSE  <= "10";
            elsif rx_error_cnt_ovf_i = '1' then
               LOST_CAUSE  <= "01";
            elsif NO_SIGNAL = '1' then
               LOST_CAUSE  <= "00";
            end if;

         end if;
      end if;
   end process p_comb_state;

--#######################################################################################--
--------------------------------------- RX processes --------------------------------------
--#######################################################################################--

-------------------------------------------------------------------------------------------
   -- RX words receive counter process
   p_rx_words_counter : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         rx_words_cnt   <= (others => '0');
         rx_new_word_r  <= '0';
      elsif rising_edge(CLK) then
         rx_new_word_r  <= RX_NEW_WORD;

         if ((RX_NEW_WORD = '1' and rx_new_word_r = '0' ) or RX_NEW_WORD = '1' ) and rx_words_cnt < C_MAX_RX_WORDS then    -- when a new word is received and lower than 16384 words receive
            rx_words_cnt <= rx_words_cnt + 1;                                                   -- Increment RX words counter by 1
         else
            rx_words_cnt <= (others => '0');                                                    -- else reset RX words counter
         end if;

      end if;
   end process p_rx_words_counter;


-------------------------------------------------------------------------------------------
   --! RX error counter process
   p_rxerr_counter : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         rx_error_cnt_i          <= (others => '0');
         rx_error_cnt_ovf_i      <= '0';
         detected_rxerr_word_r   <= '0';

      elsif rising_edge(CLK) then

         detected_rxerr_word_r   <= DETECTED_RXERR_WORD;

         if LANE_RESET = '1' or LANE_RESET_DL = '1' or current_state = CONNECTED_ST then -- Reset RXERR word counter to 0
            rx_error_cnt_i       <= (others => '0');
            rx_error_cnt_ovf_i   <= '0';

         elsif current_state = ACTIVE_ST then

            -- When 16384 words are received and a single RXERR control word is detected on 32-bit data
            if rx_words_cnt = C_MAX_RX_WORDS and ((DETECTED_RXERR_WORD = '1' and detected_rxerr_word_r = '0') or DETECTED_RXERR_WORD = '1')then
               rx_error_cnt_i <= rx_error_cnt_i;         -- do not increment RXERR word counter (counter = +1-1)
            -- When 16384 words are received and a single RXERR control word is detected on 32-bit data
            elsif rx_words_cnt = C_MAX_RX_WORDS and rx_error_cnt_i /= x"00" then
               rx_error_cnt_i <= rx_error_cnt_i - 1;         -- do not increment RXERR word counter (counter = +1-1)
            -- When a RXERR control word is detected on 32-bit data
            elsif rx_words_cnt <= C_MAX_RX_WORDS and ((DETECTED_RXERR_WORD = '1' and detected_rxerr_word_r = '0') or DETECTED_RXERR_WORD = '1') then
               if rx_error_cnt_i = C_MAX_RXERR_CTRL_WORDS then    -- Overflow gestion
                  rx_error_cnt_ovf_i   <= '1';
                  rx_error_cnt_i       <= (others => '1');        -- Lock to the max value 0xFF
               else
                  rx_error_cnt_ovf_i   <= '0';
                  rx_error_cnt_i       <= rx_error_cnt_i + 1;     -- increment RXERR word counter to 1
               end if;
            end if;
         end if;

      end if;
   end process p_rxerr_counter;

-------------------------------------------------------------------------------------------
   -- init_timeout_counter process
   p_init_timeout_counter : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         init_timeout_cnt     <= (others => '0');
         init_timeout_reaches <= '0';
      elsif rising_edge(CLK) then

         if enable_init_cnt = '1' then                      -- When the initialisation timeout counter is launched (In STARTED_ST)
            if init_timeout_cnt >= C_32US_AT_150MHZ then    -- When counter reaches 32us (time to send 5000 words with 5Gbits/s)
               init_timeout_reaches <= '1';
            else
               init_timeout_cnt  <= init_timeout_cnt+1;     -- increment counter
            end if;
         else                                               -- When the initialisation timeout counter is reseted (In ACTIVE_ST and CLEAR_LINE_ST)
            init_timeout_cnt     <= (others => '0');        -- reset counter
            init_timeout_reaches <= '0';                    -- Reset flag timeout
         end if;

      end if;
   end process p_init_timeout_counter;

-------------------------------------------------------------------------------------------
   -- Detection 3 consecutive LOST_SIGNAL process
   p_loss_signal_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         lost_signal_x3       <= '0';
         loss_signal_x3_cnt   <= "00";
      elsif rising_edge(CLK) then

         -- if the current_state signal is stable and the FSM is in ACTIVE_ST or LOSS_OF_SIGNAL_ST or PREPARE_STANDBY_ST state
         if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = LOSS_OF_SIGNAL_ST or current_state = PREPARE_STANDBY_ST) then

            if (RX_NEW_WORD = '1' and rx_new_word_r = '0')  or RX_NEW_WORD = '1' then        -- when a new word is received
               if DETECTED_LOSS_SIGNAL = '1' then                      -- and a LOSS_SIGNAL word is detected
                  if loss_signal_x3_cnt = "01" then                    -- and the cnt value is equal to 2
                     lost_signal_x3       <= '1';                      -- the transition condition is set to '1'
                     loss_signal_x3_cnt   <= "00";                     -- and the counter is set to 0
                  else
                     lost_signal_x3       <= '0';                      -- else the transition condition is set to '0'
                     loss_signal_x3_cnt   <= loss_signal_x3_cnt+1;     -- and the counter is incremented by 1
                  end if;
               else
                  lost_signal_x3          <= '0';                      -- when LOSS_SIGNAL word not detected trasition condition set to '0'
                  loss_signal_x3_cnt      <= "00";                     -- and the counter is set to 0
               end if;
            end if;
         else
            lost_signal_x3       <= '0';                               -- When a transition state is detected or the FSM is not in the right state transition condition is set to '0'
            loss_signal_x3_cnt   <= "00";                              -- and the counter is set to 0
         end if;
      end if;
   end process p_loss_signal_detection;

-------------------------------------------------------------------------------------------
   -- Detection 3 consecutive STANDBY process
   p_standby_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         standby_signal_x3       <= '0';
         standby_signal_x3_cnt   <= "00";
      elsif rising_edge(CLK) then

         -- if the current_state signal is stable and the FSM is in ACTIVE_ST or LOSS_OF_SIGNAL_ST or PREPARE_STANDBY_ST state
         if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = LOSS_OF_SIGNAL_ST or current_state = PREPARE_STANDBY_ST) then

            if (RX_NEW_WORD = '1' and rx_new_word_r = '0')  or RX_NEW_WORD = '1' then             -- when a new word is received
               if DETECTED_STANDBY = '1' then                               -- and a STANDBY word is detected
                  if standby_signal_x3_cnt = "01" then                      -- and the cnt value is equal to 2
                     standby_signal_x3       <= '1';                        -- the transition condition is set to '1'
                     standby_signal_x3_cnt   <= "00";                       -- and the counter is set to 0
                  else
                     standby_signal_x3       <= '0';                        -- else the transition condition is set to '0'
                     standby_signal_x3_cnt   <= standby_signal_x3_cnt+1;    -- and the counter is incremented by 1
                  end if;
               else
                  standby_signal_x3          <= '0';                        -- when STANDBY word not detected trasition condition set to '0'
                  standby_signal_x3_cnt      <= "00";                       -- and the counter is set to 0
               end if;
            end if;
         else
            standby_signal_x3       <= '0';                                 -- When a transition state is detected or the FSM is not in the right state transition condition is set to '0'
            standby_signal_x3_cnt   <= "00";                                -- and the counter is set to 0
         end if;
      end if;
   end process p_standby_detection;

-------------------------------------------------------------------------------------------
   -- INIT1 detection process
   p_init1_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         init1_rxed           <= '0';
         init1_rxed_r        <= '0';
         inv_init1_rxed_x3    <= '0';
         detected_init1_r     <= '0';
         detected_inv_init1_r <= '0';
         inv_init1_rxed_cnt   <= "00";
      elsif rising_edge(CLK) then
         detected_init1_r     <= DETECTED_INIT1;
         detected_inv_init1_r <= DETECTED_INV_INIT1;
         init1_rxed_r         <= init1_rxed;

         -- States for detection of at least one INIT1 is received and no rx error is detected
         if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) and DETECTED_RXERR_WORD = '0' then

            if (DETECTED_INV_INIT1 = '1' and detected_inv_init1_r = '0') or DETECTED_INV_INIT1 = '1' then   -- INIT1 inversed detection condition
               if inv_init1_rxed_cnt >= "10" then                             -- and the counter reaches 3
                  inv_init1_rxed_cnt <= "00";                                 -- reset counter
                  inv_init1_rxed_x3  <= '1';                                  -- Set to '1' the transition condition to INVERT_RX_POLARITY_ST
               else
                  inv_init1_rxed_cnt <= inv_init1_rxed_cnt+1;                 -- else increment counter by 1
                  inv_init1_rxed_x3  <= '0';                                  -- Set to '0' the transition condition to INVERT_RX_POLARITY_ST
               end if;
            end if;

            if (DETECTED_INIT1 = '1' and detected_init1_r = '0' ) or DETECTED_INIT1 = '1' then           -- INIT1 detection condition
               init1_rxed  <= '1';                                            -- Set to '1' transition condition to CONNECTING_ST or LOSS_OF_SIGNAL_ST
            end if;
         else
            init1_rxed           <= '0';                                      -- else reset flags and counter
            inv_init1_rxed_cnt   <= "00";
            inv_init1_rxed_x3    <= '0';
         end if;
      end if;
   end process p_init1_detection;

-------------------------------------------------------------------------------------------
   -- INIT2 detection process
   p_init2_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         inv_init2_rxed_x3    <= '0';
         inv_init2_rxed_cnt   <= "00";
         init2_rxed_cnt       <= "00";
         init2_rxed_x3        <= '0';
         detected_inv_init2_r <= '0';
         detected_init2_r     <= '0';
         init2_rxed           <= '0';
      elsif rising_edge(CLK) then
         detected_init2_r     <= DETECTED_INIT2;
         detected_inv_init2_r <= DETECTED_INV_INIT2;

         -- States for detection of at least one INIT2 is received and no rx error is detected
         if current_state = current_state_r and (current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST or current_state = CONNECTING_ST) and DETECTED_RXERR_WORD = '0' then

            if (DETECTED_INV_INIT2 = '1' and detected_inv_init2_r = '0') or DETECTED_INV_INIT2 = '1' then   -- INIT2 inversed detection condition
               if inv_init2_rxed_cnt >= "10" then                             -- and the counter reaches 3
                  inv_init2_rxed_cnt   <= "00";                               -- reset counter
                  inv_init2_rxed_x3    <= '1';                                -- Set to '1' the transition condition to INVERT_RX_POLARITY_ST
               else
                  inv_init2_rxed_cnt   <= inv_init2_rxed_cnt+1;               -- else increment by 1
                  inv_init2_rxed_x3    <= '0';                                -- Set to '0' the transition condition to INVERT_RX_POLARITY_ST
               end if;
            end if;

            if (DETECTED_INIT2 = '1' and detected_init2_r = '0') or DETECTED_INIT2 = '1' then           -- INIT2 detection condition
               init2_rxed  <= '1';
               if init2_rxed_cnt >= "10" then                                 -- and the counter reaches 3
                  init2_rxed_cnt <= "00";                                     -- reset counter
                  init2_rxed_x3  <= '1';                                      -- Set to '1' the transition condition to CONNECTING_ST
               else
                  init2_rxed_cnt <= init2_rxed_cnt+1;                         -- else increment counter by 1
                  init2_rxed_x3  <= '0';                                      -- Set to '0' the transition condition to CONNECTING_ST
               end if;
            end if;

         else
            inv_init2_rxed_x3    <= '0';                                      -- else reset flags and counters
            inv_init2_rxed_cnt   <= "00";
            init2_rxed_cnt       <= "00";
            init2_rxed_x3        <= '0';
            init2_rxed           <= '0';
         end if;
      end if;
   end process p_init2_detection;

-------------------------------------------------------------------------------------------
   -- INIT3 detection process
   p_init3_detection : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         init3_rxed_x3    <= '0';
         init3_rxed_cnt   <= "00";
         detected_init3_r <= '0';
         comma_k287_rxed_r <= '0';
      elsif rising_edge(CLK) then
         detected_init3_r  <= DETECTED_INIT3;
         comma_k287_rxed_r <= COMMA_K287_RXED;

         -- States for detection of INIT3 is received and no rx error is detected
         if current_state = current_state_r and (current_state = CONNECTING_ST or current_state = CONNECTED_ST) and DETECTED_RXERR_WORD = '0' then

            if (DETECTED_INIT3 = '1' and detected_init3_r = '0') or DETECTED_INIT3 = '1' then  -- INIT3 detection condition
               if init3_rxed_cnt = "10" then                         -- and counter reaches 3
                  init3_rxed_cnt   <= "00";                          -- reset counter
                  init3_rxed_x3    <= '1';                           -- Set to '1' transition condition to CONNECTING_ST or ACTIVE_ST
               else
                  init3_rxed_cnt   <= init3_rxed_cnt+1;              -- else increment counter by 1
                  init3_rxed_x3    <= '0';                           -- Set to '0' transition condition to CONNECTING_ST or ACTIVE_ST
               end if;
            end if;
         else
            init3_rxed_cnt   <= "00";                                -- reset flag and counter
            init3_rxed_x3    <= '0';
         end if;

      end if;
   end process p_init3_detection;

-------------------------------------------------------------------------------------------
   -- Process for detection the reception of 1023 words including the reception of at least on INIT1 or INIT2 without RXERR control words
   p_init1_or_init2_detection_without_rx_error : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         rxed_1023_word       <= '0';
         rxed_1023_word_cnt   <= (others => '0');

      elsif rising_edge(CLK) then

         -- if the current_state signal is stable and the FSM is in STARTED_ST or INVERT_ST state
         if current_state = current_state_r and (current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then

            if ((RX_NEW_WORD = '1' and rx_new_word_r = '0') or RX_NEW_WORD = '1') then            -- when new word is received
               if DETECTED_RXERR_WORD = '0' then                           -- and no error has occurred
                  if rxed_1023_word_cnt >= C_1023_WORDS-1 then             -- when 1023 words are receive without error
                     if init1_rxed = '1' or init2_rxed = '1'  then         -- when at least one INIT1 or INIT2 is received and no RXERR detected
                        rxed_1023_word    <= '1';                          -- set transition condition to '1'
                     else
                        rxed_1023_word    <= '0';                          -- set transition condition to '0'
                     end if;
                  else
                     rxed_1023_word_cnt   <= rxed_1023_word_cnt+1;         -- increment counter by 1
                     rxed_1023_word       <= '0';                          -- set transition condition to '0'
                  end if;
               else
                  rxed_1023_word_cnt      <= (others => '0');              -- reset counter
                  rxed_1023_word          <= '0';
               end if;
            end if;
         else
            rxed_1023_word_cnt   <= (others => '0');                       -- reset counter
            rxed_1023_word       <= '0';                                   -- set transition condition to '0'
         end if;
      end if;
   end process p_init1_or_init2_detection_without_rx_error;

-------------------------------------------------------------------------------------------
   -- RXERR word send to data_link when FSM leave ACTIVE_ST process
   p_send_rx_error_word : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         SEND_RXERR  <= '0';
      elsif rising_edge(CLK) then
         if current_state /= ACTIVE_ST and current_state_r = ACTIVE_ST then   -- when the FSM get out from the ACTIVE_ST
            SEND_RXERR  <= '1';                                               -- Set flag to '1' in order to send RXERR control word to Data-link layer
         else
            SEND_RXERR  <= '0';                                               -- else set flag to '0'
         end if;
      end if;
   end process p_send_rx_error_word;


-- Outputs
CDR            <= cdr_i;
RX_ERROR_CNT   <= std_logic_vector(rx_error_cnt_i);
RX_ERROR_OVF   <= rx_error_cnt_ovf_i;

end architecture rtl;
