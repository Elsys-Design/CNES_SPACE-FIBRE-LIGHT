LIBRARY ieee ;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--library work;

entity tb_lane_init_fsm is
end entity;

architecture tb of tb_lane_init_fsm is

component lane_init_fsm is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP
      -- FROM/TO Data-link layer
      LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer.

      -- RX signals
      NO_SIGNAL                        : in  std_logic;                       --! Flag no signal are received
      RX_NEW_WORD                      : in  std_logic;                       --! Flag new word has been received
      DETECTED_INIT1                   : in  std_logic;                       --! Flag INIT1 control word rxed
      DETECTED_INIT2                   : in  std_logic;                       --! Flag INIT2 control word rxed
      DETECTED_INIT3                   : in  std_logic;                       --! Flag INIT3 control word rxed
      DETECTED_INV_INIT1               : in  std_logic;                       --! Flag INV_INIT1 control word rxed
      DETECTED_INV_INIT2               : in  std_logic;                       --! Flag INV_INIT2 control word rxed
      DETECTED_RXERR_WORD              : in  std_logic;                       --! Flag RXERR detected
      DETECTED_LOSS_SIGNAL             : in  std_logic;                       --! Flag LOSS_SINGAL control word detected
      DETECTED_STANDBY                 : in  std_logic;                       --! Flag STANDBY control word detected
      COMMA_K287_RXED                  : in  std_logic;                       --! Flag Comma K28.7 has been received
      RECEIVER_DISABLED                : out std_logic;                       --! flag to enabled RX function of HSSL IP
      CDR                              : out std_logic;                       --! Flag to enabled CDR function of HSSL IP
      SEND_RXERR                       : out std_logic;                       --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
      INVERT_RX_BITS                   : out std_logic;                       --! Flag to Invert rx bit received
      NO_SIGNAL_DETECTION_ENABLED      : out std_logic;                       --! Flag to enable the no signal function

      -- TX signals
      STANDBY_SIGNAL_X32               : in  std_logic;                       --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32                  : in  std_logic;                       --! Flag LOST_SIGNAL control word has been send x32
      TRANSMITTER_DISABLED             : out std_logic;                       --! flag to enabled TX fonction of HSSL IP
      SEND_INIT1_CTRL_WORD             : out std_logic;                       --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD             : out std_logic;                       --! Flag to send control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD             : out std_logic;                       --! Flag to send control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA               : out std_logic;                       --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS       : out std_logic;                       --! Flag to send STANDBY control word x32
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   : out std_logic;                       --! Flag to send LOSS_SIGNAL control word x32
      LOST_CAUSE                       : out std_logic_vector(01 downto 00);  --! Flag to indicate the reason of the LOST_SIGNAL

      -- PARAMETERS and STATUS
      LANE_START                       : in  std_logic;                       --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                       --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                       --! Asserts or de-asserts LaneReset for the lane
      LANE_STATE                       : out std_logic_vector(03 downto 00);  --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic                        --! Overflow flag of the RX_ERROR_CNT
   );
end component;


----------------------------- Stimulus signals
constant periode                       : time := 6.667 ns;
----- inputs
signal RST_N                           : std_logic := '1';
signal CLK                             : std_logic := '0';
signal LANE_RESET_DL                   : std_logic := '0';
------ RX signals
signal NO_SIGNAL                       : std_logic := '1';
signal RX_NEW_WORD                     : std_logic := '0';
signal DETECTED_INIT1                  : std_logic := '0';
signal DETECTED_INIT2                  : std_logic := '0';
signal DETECTED_INIT3                  : std_logic := '0';
signal DETECTED_INV_INIT1              : std_logic := '0';
signal DETECTED_INV_INIT2              : std_logic := '0';
signal DETECTED_RXERR_WORD             : std_logic := '0';
signal DETECTED_LOSS_SIGNAL            : std_logic := '0';
signal DETECTED_STANDBY                : std_logic := '0';
signal COMMA_K287_RXED                 : std_logic := '0';
   ------ TX signals
signal STANDBY_SIGNAL_X32              : std_logic := '0';
signal LOST_SIGNAL_X32                 : std_logic := '0';
   ------ PARAMETERS
signal LANE_START                      : std_logic := '0';
signal AUTOSTART                       : std_logic := '0';
signal LANE_RESET                      : std_logic := '0';

----- Outputs
   ------ RX signals
signal RECEIVER_DISABLED                : std_logic := '0';
signal CDR                             : std_logic := '0';
signal SEND_RXERR                      : std_logic := '0';
signal INVERT_RX_BITS                  : std_logic := '0';
signal NO_SIGNAL_DETECTION_ENABLED     : std_logic := '0';
   ------ TX signals
signal TRANSMITTER_DISABLED             : std_logic := '0';
signal SEND_INIT1_CTRL_WORD            : std_logic := '0';
signal SEND_INIT2_CTRL_WORD            : std_logic := '0';
signal SEND_INIT3_CTRL_WORD            : std_logic := '0';
signal ENABLE_TRANSM_DATA              : std_logic := '0';
signal SEND_32_STANDBY_CTRL_WORDS      : std_logic := '0';
signal SEND_32_LOSS_SIGNAL_CTRL_WORDS  : std_logic := '0';
signal LOST_CAUSE                      : std_logic_vector(01 downto 00);
   ------ STATUS
signal LANE_STATE                      : std_logic_vector(03 downto 00) := x"0";
signal RX_ERROR_CNT                    : std_logic_vector(07 downto 00) := x"00";
signal RX_ERROR_OVF                    : std_logic := '0';

begin

DUT : lane_init_fsm
   port map(
      RST_N                            => RST_N,
      CLK                              => CLK,
      -- FROM/TO Data-link layer
      LANE_RESET_DL                    => LANE_RESET_DL,
      -- RX signals
      NO_SIGNAL                        => NO_SIGNAL,
      RX_NEW_WORD                      => RX_NEW_WORD,
      DETECTED_INIT1                   => DETECTED_INIT1,
      DETECTED_INIT2                   => DETECTED_INIT2,
      DETECTED_INIT3                   => DETECTED_INIT3,
      DETECTED_INV_INIT1               => DETECTED_INV_INIT1,
      DETECTED_INV_INIT2               => DETECTED_INV_INIT2,
      DETECTED_RXERR_WORD              => DETECTED_RXERR_WORD,
      DETECTED_LOSS_SIGNAL             => DETECTED_LOSS_SIGNAL,
      DETECTED_STANDBY                 => DETECTED_STANDBY,
      COMMA_K287_RXED                  => COMMA_K287_RXED,
      RECEIVER_DISABLED                 => RECEIVER_DISABLED,
      CDR                              => CDR,
      SEND_RXERR                       => SEND_RXERR,
      INVERT_RX_BITS                   => INVERT_RX_BITS,
      NO_SIGNAL_DETECTION_ENABLED      => NO_SIGNAL_DETECTION_ENABLED,
      -- TX signals
      STANDBY_SIGNAL_X32               => STANDBY_SIGNAL_X32,
      LOST_SIGNAL_X32                  => LOST_SIGNAL_X32,
      TRANSMITTER_DISABLED              => TRANSMITTER_DISABLED,
      SEND_INIT1_CTRL_WORD             => SEND_INIT1_CTRL_WORD,
      SEND_INIT2_CTRL_WORD             => SEND_INIT2_CTRL_WORD,
      SEND_INIT3_CTRL_WORD             => SEND_INIT3_CTRL_WORD,
      ENABLE_TRANSM_DATA               => ENABLE_TRANSM_DATA,
      SEND_32_STANDBY_CTRL_WORDS       => SEND_32_STANDBY_CTRL_WORDS,
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   => SEND_32_LOSS_SIGNAL_CTRL_WORDS,
      LOST_CAUSE                       => LOST_CAUSE,
      -- PARAMETERS and STATUS
      LANE_START                       => LANE_START,
      AUTOSTART                        => AUTOSTART,
      LANE_RESET                       => LANE_RESET,
      LANE_STATE                       => LANE_STATE,
      RX_ERROR_CNT                     => RX_ERROR_CNT,
      RX_ERROR_OVF                     => RX_ERROR_OVF);


-- generate clock 150 MHz
horloge : process
begin
   CLK   <= not CLK;
   wait for periode/2;
end process;

scenario : process
begin
-- LANE_START
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 20 us;
   AUTOSTART  <= '1';
   
   wait for 20 ns;
   NO_SIGNAL   <= '0';
   
   -- STARTED_ST to INVERT_ST
   wait until rising_edge(CLK);
   test_loop : for k in 0 to 2 loop
      RX_NEW_WORD    <= '1';
      DETECTED_INV_INIT1 <= '1';
      wait until rising_edge(CLK);
      RX_NEW_WORD    <= '0';
      DETECTED_INV_INIT1 <= '0';
      wait until rising_edge(CLK);
   end loop;
   
   wait until rising_edge(CLK);
   
   -- INVERT_ST to CONNECTING_ST
   test1_loop : for k in 0 to 1022 loop
      RX_NEW_WORD    <= '1';
      DETECTED_INIT1 <= '1';
      wait until rising_edge(CLK);
      RX_NEW_WORD    <= '0';
      DETECTED_INIT1 <= '0';
      wait until rising_edge(CLK);
   end loop;
   
   wait until rising_edge(CLK);
   
   -- CONNECTING_ST to CONNECTED_ST
   test2_loop : for k in 0 to 2 loop
      RX_NEW_WORD    <= '1';
      DETECTED_INIT2 <= '1';
      wait until rising_edge(CLK);
      RX_NEW_WORD    <= '0';
      DETECTED_INIT2 <= '0';
      wait until rising_edge(CLK);
   end loop;
   
   wait until rising_edge(CLK);
   
   -- CONNECTED_ST to ACTIVE_ST
   test3_loop : for k in 0 to 2 loop
      RX_NEW_WORD    <= '1';
      DETECTED_INIT3 <= '1';
      wait until rising_edge(CLK);
      RX_NEW_WORD    <= '0';
      DETECTED_INIT3 <= '0';
      wait until rising_edge(CLK);
   end loop;
   
   wait for 10 us;
   
   
   AUTOSTART   <= '0';
   -- In ACTIVE_ST compteur RXERR
   -- test4_loop : for k in 0 to 256 loop
      -- RX_NEW_WORD    <= '1';
      -- DETECTED_RXERR_WORD <= '1';
      -- wait until rising_edge(CLK);
      -- RX_NEW_WORD    <= '0';
      -- DETECTED_RXERR_WORD <= '0';
      -- wait until rising_edge(CLK);
   -- end loop;
   
   -- wait until rising_edge(CLK);
   
   wait;   
end process;

end tb;