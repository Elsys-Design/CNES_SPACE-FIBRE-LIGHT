// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC_NPS4_DEFINES_VH
`else
`define B_NOC_NPS4_DEFINES_VH

// Look-up table parameters
//

`define NOC_NPS4_ADDR_N  37
`define NOC_NPS4_ADDR_SZ 32
`define NOC_NPS4_DATA_SZ 32

// Attribute addresses
//

`define NOC_NPS4__REG_DST_ID_P0    32'h00000000
`define NOC_NPS4__REG_DST_ID_P0_SZ 12

`define NOC_NPS4__REG_DST_ID_P1    32'h00000001
`define NOC_NPS4__REG_DST_ID_P1_SZ 12

`define NOC_NPS4__REG_DST_ID_P2    32'h00000002
`define NOC_NPS4__REG_DST_ID_P2_SZ 12

`define NOC_NPS4__REG_DST_ID_P3    32'h00000003
`define NOC_NPS4__REG_DST_ID_P3_SZ 12

`define NOC_NPS4__REG_HBM2NOC_P0_P0_VCA_TOKEN    32'h00000004
`define NOC_NPS4__REG_HBM2NOC_P0_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P0_P1_VCA_TOKEN    32'h00000005
`define NOC_NPS4__REG_HBM2NOC_P0_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P0_P2_VCA_TOKEN    32'h00000006
`define NOC_NPS4__REG_HBM2NOC_P0_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P0_P3_VCA_TOKEN    32'h00000007
`define NOC_NPS4__REG_HBM2NOC_P0_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P1_P0_VCA_TOKEN    32'h00000008
`define NOC_NPS4__REG_HBM2NOC_P1_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P1_P1_VCA_TOKEN    32'h00000009
`define NOC_NPS4__REG_HBM2NOC_P1_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P1_P2_VCA_TOKEN    32'h0000000a
`define NOC_NPS4__REG_HBM2NOC_P1_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P1_P3_VCA_TOKEN    32'h0000000b
`define NOC_NPS4__REG_HBM2NOC_P1_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P2_P0_VCA_TOKEN    32'h0000000c
`define NOC_NPS4__REG_HBM2NOC_P2_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P2_P1_VCA_TOKEN    32'h0000000d
`define NOC_NPS4__REG_HBM2NOC_P2_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P2_P2_VCA_TOKEN    32'h0000000e
`define NOC_NPS4__REG_HBM2NOC_P2_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P2_P3_VCA_TOKEN    32'h0000000f
`define NOC_NPS4__REG_HBM2NOC_P2_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P3_P0_VCA_TOKEN    32'h00000010
`define NOC_NPS4__REG_HBM2NOC_P3_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P3_P1_VCA_TOKEN    32'h00000011
`define NOC_NPS4__REG_HBM2NOC_P3_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P3_P2_VCA_TOKEN    32'h00000012
`define NOC_NPS4__REG_HBM2NOC_P3_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_HBM2NOC_P3_P3_VCA_TOKEN    32'h00000013
`define NOC_NPS4__REG_HBM2NOC_P3_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P0_P0_VCA_TOKEN    32'h00000014
`define NOC_NPS4__REG_NOC2HBM_P0_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P0_P1_VCA_TOKEN    32'h00000015
`define NOC_NPS4__REG_NOC2HBM_P0_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P0_P2_VCA_TOKEN    32'h00000016
`define NOC_NPS4__REG_NOC2HBM_P0_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P0_P3_VCA_TOKEN    32'h00000017
`define NOC_NPS4__REG_NOC2HBM_P0_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P1_P0_VCA_TOKEN    32'h00000018
`define NOC_NPS4__REG_NOC2HBM_P1_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P1_P1_VCA_TOKEN    32'h00000019
`define NOC_NPS4__REG_NOC2HBM_P1_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P1_P2_VCA_TOKEN    32'h0000001a
`define NOC_NPS4__REG_NOC2HBM_P1_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P1_P3_VCA_TOKEN    32'h0000001b
`define NOC_NPS4__REG_NOC2HBM_P1_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P2_P0_VCA_TOKEN    32'h0000001c
`define NOC_NPS4__REG_NOC2HBM_P2_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P2_P1_VCA_TOKEN    32'h0000001d
`define NOC_NPS4__REG_NOC2HBM_P2_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P2_P2_VCA_TOKEN    32'h0000001e
`define NOC_NPS4__REG_NOC2HBM_P2_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P2_P3_VCA_TOKEN    32'h0000001f
`define NOC_NPS4__REG_NOC2HBM_P2_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P3_P0_VCA_TOKEN    32'h00000020
`define NOC_NPS4__REG_NOC2HBM_P3_P0_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P3_P1_VCA_TOKEN    32'h00000021
`define NOC_NPS4__REG_NOC2HBM_P3_P1_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P3_P2_VCA_TOKEN    32'h00000022
`define NOC_NPS4__REG_NOC2HBM_P3_P2_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC2HBM_P3_P3_VCA_TOKEN    32'h00000023
`define NOC_NPS4__REG_NOC2HBM_P3_P3_VCA_TOKEN_SZ 32

`define NOC_NPS4__REG_NOC_CTL    32'h00000024
`define NOC_NPS4__REG_NOC_CTL_SZ 1

`endif  // B_NOC_NPS4_DEFINES_VH