-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 18/06/2025
--
-- Description : This module allows realigning the beginnings of words so
--               that they start on byte 0 or 4.
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.all;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_word_alignment is
   port (
      RST_N                            : in  std_logic;                                           --! global reset
      CLK                              : in  std_logic;                                           --! Clock generated by HSSL IP
      -- TO lane_ctrl_word_detection
      DATA_RX_TO_LCWD                  : out std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! 64-bit data to lane_ctrl_word_detect
      VALID_K_CHARAC_TO_LCWD            : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! 8-bit valid K character flags to lane_ctrl_word_detect
      DATA_RDY_TO_LCWD                 : out std_logic;                                           --! Data valid flag to lane_ctrl_word_detect
      -- FROM MANUFACTURER IP
      DATA_RX_FROM_IP                  : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! 64-bit data from HSSL IP
      VALID_K_CHARAC_FROM_IP            : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! 8-bit valid K character flags from HSSL IP
      RX_WORD_IS_ALIGNED_FROM_IP       : in  std_logic;                                           --! RX word is aligned from HSSL IP
      COMMA_DET_FROM_IP                : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0)   --! Flag indicates that a comma is detected on the word receive
   );
end ppl_64_word_alignment;

architecture rtl of ppl_64_word_alignment is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------

  signal reg_data       : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal reg_k_char     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal alignment_byte : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_rx_realignment
-- Description: Align the words so that they are at the beginning of the bus.
---------------------------------------------------------
  p_rx_realignment: process(CLK,RST_N)
  begin
    if RST_N = '0' then
      DATA_RX_TO_LCWD        <= (others => '0');
      VALID_K_CHARAC_TO_LCWD  <= (others => '0');
      DATA_RDY_TO_LCWD       <= '0';
      alignment_byte         <= (others => '0');
      reg_data               <= (others => '0');
      reg_k_char             <= (others => '0');
    elsif rising_edge(CLK) then
      if RX_WORD_IS_ALIGNED_FROM_IP ='1' then
        if alignment_byte(7) = '1' or (COMMA_DET_FROM_IP(7) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "10000000";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(7*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 7*8)  ;
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(7-1 downto 0) & reg_k_char(7);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(6) = '1' or (COMMA_DET_FROM_IP(6) = '1' and alignment_byte= std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "01000000";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(6*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 6*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(6-1 downto 0) & reg_k_char(7 downto 6);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(5) = '1' or (COMMA_DET_FROM_IP(5) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00100000";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(5*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 5*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(5-1 downto 0) & reg_k_char(7 downto 5);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(4) = '1' or (COMMA_DET_FROM_IP(4) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00010000";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(4*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 4*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(4-1 downto 0) & reg_k_char(7 downto 4);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(3) = '1' or (COMMA_DET_FROM_IP(3) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00001000";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(3*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 3*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(3-1 downto 0) & reg_k_char(7 downto 3);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(2) = '1' or (COMMA_DET_FROM_IP(2) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00000100";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(2*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 2*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(2-1 downto 0) & reg_k_char(7 downto 2);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(1) = '1' or (COMMA_DET_FROM_IP(1) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00000010";
          reg_data                                       <= DATA_RX_FROM_IP;
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP(1*8-1 downto 0) & reg_data(C_BYTE_BY_WORD_LENGTH*8-1 downto 1*8);
          reg_k_char                                     <= VALID_K_CHARAC_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP(1-1 downto 0) & reg_k_char(7 downto 1);
          DATA_RDY_TO_LCWD                               <= '1';
        elsif alignment_byte(0) = '1' or (COMMA_DET_FROM_IP(0) = '1' and alignment_byte = std_logic_vector(to_unsigned(0,alignment_byte'length)))  then
          alignment_byte                                 <= "00000001";
          DATA_RX_TO_LCWD                                <= DATA_RX_FROM_IP;
          VALID_K_CHARAC_TO_LCWD                          <= VALID_K_CHARAC_FROM_IP;
          DATA_RDY_TO_LCWD                               <= '1';
        end if;
      else
        DATA_RX_TO_LCWD        <= (others => '0');
        VALID_K_CHARAC_TO_LCWD  <= (others => '0');
        DATA_RDY_TO_LCWD       <= '0';
        alignment_byte         <= (others => '0');
        reg_data               <= (others => '0');
        reg_k_char             <= (others => '0');
      end if;
    end if;
  end process p_rx_realignment;
  
end architecture rtl;