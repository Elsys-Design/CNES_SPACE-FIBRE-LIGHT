// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_CMACE4_DEFINES_VH
`else
`define B_CMACE4_DEFINES_VH

// Look-up table parameters
//

`define CMACE4_ADDR_N  84
`define CMACE4_ADDR_SZ 32
`define CMACE4_DATA_SZ 152

// Attribute addresses
//

`define CMACE4__CTL_PTP_TRANSPCLK_MODE    32'h00000000
`define CMACE4__CTL_PTP_TRANSPCLK_MODE_SZ 40

`define CMACE4__CTL_RX_CHECK_ACK    32'h00000001
`define CMACE4__CTL_RX_CHECK_ACK_SZ 40

`define CMACE4__CTL_RX_CHECK_PREAMBLE    32'h00000002
`define CMACE4__CTL_RX_CHECK_PREAMBLE_SZ 40

`define CMACE4__CTL_RX_CHECK_SFD    32'h00000003
`define CMACE4__CTL_RX_CHECK_SFD_SZ 40

`define CMACE4__CTL_RX_DELETE_FCS    32'h00000004
`define CMACE4__CTL_RX_DELETE_FCS_SZ 40

`define CMACE4__CTL_RX_ETYPE_GCP    32'h00000005
`define CMACE4__CTL_RX_ETYPE_GCP_SZ 16

`define CMACE4__CTL_RX_ETYPE_GPP    32'h00000006
`define CMACE4__CTL_RX_ETYPE_GPP_SZ 16

`define CMACE4__CTL_RX_ETYPE_PCP    32'h00000007
`define CMACE4__CTL_RX_ETYPE_PCP_SZ 16

`define CMACE4__CTL_RX_ETYPE_PPP    32'h00000008
`define CMACE4__CTL_RX_ETYPE_PPP_SZ 16

`define CMACE4__CTL_RX_FORWARD_CONTROL    32'h00000009
`define CMACE4__CTL_RX_FORWARD_CONTROL_SZ 40

`define CMACE4__CTL_RX_IGNORE_FCS    32'h0000000a
`define CMACE4__CTL_RX_IGNORE_FCS_SZ 40

`define CMACE4__CTL_RX_MAX_PACKET_LEN    32'h0000000b
`define CMACE4__CTL_RX_MAX_PACKET_LEN_SZ 15

`define CMACE4__CTL_RX_MIN_PACKET_LEN    32'h0000000c
`define CMACE4__CTL_RX_MIN_PACKET_LEN_SZ 8

`define CMACE4__CTL_RX_OPCODE_GPP    32'h0000000d
`define CMACE4__CTL_RX_OPCODE_GPP_SZ 16

`define CMACE4__CTL_RX_OPCODE_MAX_GCP    32'h0000000e
`define CMACE4__CTL_RX_OPCODE_MAX_GCP_SZ 16

`define CMACE4__CTL_RX_OPCODE_MAX_PCP    32'h0000000f
`define CMACE4__CTL_RX_OPCODE_MAX_PCP_SZ 16

`define CMACE4__CTL_RX_OPCODE_MIN_GCP    32'h00000010
`define CMACE4__CTL_RX_OPCODE_MIN_GCP_SZ 16

`define CMACE4__CTL_RX_OPCODE_MIN_PCP    32'h00000011
`define CMACE4__CTL_RX_OPCODE_MIN_PCP_SZ 16

`define CMACE4__CTL_RX_OPCODE_PPP    32'h00000012
`define CMACE4__CTL_RX_OPCODE_PPP_SZ 16

`define CMACE4__CTL_RX_PAUSE_DA_MCAST    32'h00000013
`define CMACE4__CTL_RX_PAUSE_DA_MCAST_SZ 48

`define CMACE4__CTL_RX_PAUSE_DA_UCAST    32'h00000014
`define CMACE4__CTL_RX_PAUSE_DA_UCAST_SZ 48

`define CMACE4__CTL_RX_PAUSE_SA    32'h00000015
`define CMACE4__CTL_RX_PAUSE_SA_SZ 48

`define CMACE4__CTL_RX_PROCESS_LFI    32'h00000016
`define CMACE4__CTL_RX_PROCESS_LFI_SZ 40

`define CMACE4__CTL_RX_RSFEC_AM_THRESHOLD    32'h00000017
`define CMACE4__CTL_RX_RSFEC_AM_THRESHOLD_SZ 9

`define CMACE4__CTL_RX_RSFEC_FILL_ADJUST    32'h00000018
`define CMACE4__CTL_RX_RSFEC_FILL_ADJUST_SZ 2

`define CMACE4__CTL_RX_VL_LENGTH_MINUS1    32'h00000019
`define CMACE4__CTL_RX_VL_LENGTH_MINUS1_SZ 16

`define CMACE4__CTL_RX_VL_MARKER_ID0    32'h0000001a
`define CMACE4__CTL_RX_VL_MARKER_ID0_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID1    32'h0000001b
`define CMACE4__CTL_RX_VL_MARKER_ID1_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID10    32'h0000001c
`define CMACE4__CTL_RX_VL_MARKER_ID10_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID11    32'h0000001d
`define CMACE4__CTL_RX_VL_MARKER_ID11_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID12    32'h0000001e
`define CMACE4__CTL_RX_VL_MARKER_ID12_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID13    32'h0000001f
`define CMACE4__CTL_RX_VL_MARKER_ID13_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID14    32'h00000020
`define CMACE4__CTL_RX_VL_MARKER_ID14_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID15    32'h00000021
`define CMACE4__CTL_RX_VL_MARKER_ID15_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID16    32'h00000022
`define CMACE4__CTL_RX_VL_MARKER_ID16_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID17    32'h00000023
`define CMACE4__CTL_RX_VL_MARKER_ID17_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID18    32'h00000024
`define CMACE4__CTL_RX_VL_MARKER_ID18_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID19    32'h00000025
`define CMACE4__CTL_RX_VL_MARKER_ID19_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID2    32'h00000026
`define CMACE4__CTL_RX_VL_MARKER_ID2_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID3    32'h00000027
`define CMACE4__CTL_RX_VL_MARKER_ID3_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID4    32'h00000028
`define CMACE4__CTL_RX_VL_MARKER_ID4_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID5    32'h00000029
`define CMACE4__CTL_RX_VL_MARKER_ID5_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID6    32'h0000002a
`define CMACE4__CTL_RX_VL_MARKER_ID6_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID7    32'h0000002b
`define CMACE4__CTL_RX_VL_MARKER_ID7_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID8    32'h0000002c
`define CMACE4__CTL_RX_VL_MARKER_ID8_SZ 64

`define CMACE4__CTL_RX_VL_MARKER_ID9    32'h0000002d
`define CMACE4__CTL_RX_VL_MARKER_ID9_SZ 64

`define CMACE4__CTL_TEST_MODE_PIN_CHAR    32'h0000002e
`define CMACE4__CTL_TEST_MODE_PIN_CHAR_SZ 40

`define CMACE4__CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h0000002f
`define CMACE4__CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define CMACE4__CTL_TX_DA_GPP    32'h00000030
`define CMACE4__CTL_TX_DA_GPP_SZ 48

`define CMACE4__CTL_TX_DA_PPP    32'h00000031
`define CMACE4__CTL_TX_DA_PPP_SZ 48

`define CMACE4__CTL_TX_ETHERTYPE_GPP    32'h00000032
`define CMACE4__CTL_TX_ETHERTYPE_GPP_SZ 16

`define CMACE4__CTL_TX_ETHERTYPE_PPP    32'h00000033
`define CMACE4__CTL_TX_ETHERTYPE_PPP_SZ 16

`define CMACE4__CTL_TX_FCS_INS_ENABLE    32'h00000034
`define CMACE4__CTL_TX_FCS_INS_ENABLE_SZ 40

`define CMACE4__CTL_TX_IGNORE_FCS    32'h00000035
`define CMACE4__CTL_TX_IGNORE_FCS_SZ 40

`define CMACE4__CTL_TX_IPG_VALUE    32'h00000036
`define CMACE4__CTL_TX_IPG_VALUE_SZ 4

`define CMACE4__CTL_TX_OPCODE_GPP    32'h00000037
`define CMACE4__CTL_TX_OPCODE_GPP_SZ 16

`define CMACE4__CTL_TX_OPCODE_PPP    32'h00000038
`define CMACE4__CTL_TX_OPCODE_PPP_SZ 16

`define CMACE4__CTL_TX_PTP_1STEP_ENABLE    32'h00000039
`define CMACE4__CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define CMACE4__CTL_TX_PTP_LATENCY_ADJUST    32'h0000003a
`define CMACE4__CTL_TX_PTP_LATENCY_ADJUST_SZ 11

`define CMACE4__CTL_TX_SA_GPP    32'h0000003b
`define CMACE4__CTL_TX_SA_GPP_SZ 48

`define CMACE4__CTL_TX_SA_PPP    32'h0000003c
`define CMACE4__CTL_TX_SA_PPP_SZ 48

`define CMACE4__CTL_TX_VL_LENGTH_MINUS1    32'h0000003d
`define CMACE4__CTL_TX_VL_LENGTH_MINUS1_SZ 16

`define CMACE4__CTL_TX_VL_MARKER_ID0    32'h0000003e
`define CMACE4__CTL_TX_VL_MARKER_ID0_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID1    32'h0000003f
`define CMACE4__CTL_TX_VL_MARKER_ID1_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID10    32'h00000040
`define CMACE4__CTL_TX_VL_MARKER_ID10_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID11    32'h00000041
`define CMACE4__CTL_TX_VL_MARKER_ID11_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID12    32'h00000042
`define CMACE4__CTL_TX_VL_MARKER_ID12_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID13    32'h00000043
`define CMACE4__CTL_TX_VL_MARKER_ID13_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID14    32'h00000044
`define CMACE4__CTL_TX_VL_MARKER_ID14_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID15    32'h00000045
`define CMACE4__CTL_TX_VL_MARKER_ID15_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID16    32'h00000046
`define CMACE4__CTL_TX_VL_MARKER_ID16_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID17    32'h00000047
`define CMACE4__CTL_TX_VL_MARKER_ID17_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID18    32'h00000048
`define CMACE4__CTL_TX_VL_MARKER_ID18_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID19    32'h00000049
`define CMACE4__CTL_TX_VL_MARKER_ID19_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID2    32'h0000004a
`define CMACE4__CTL_TX_VL_MARKER_ID2_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID3    32'h0000004b
`define CMACE4__CTL_TX_VL_MARKER_ID3_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID4    32'h0000004c
`define CMACE4__CTL_TX_VL_MARKER_ID4_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID5    32'h0000004d
`define CMACE4__CTL_TX_VL_MARKER_ID5_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID6    32'h0000004e
`define CMACE4__CTL_TX_VL_MARKER_ID6_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID7    32'h0000004f
`define CMACE4__CTL_TX_VL_MARKER_ID7_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID8    32'h00000050
`define CMACE4__CTL_TX_VL_MARKER_ID8_SZ 64

`define CMACE4__CTL_TX_VL_MARKER_ID9    32'h00000051
`define CMACE4__CTL_TX_VL_MARKER_ID9_SZ 64

`define CMACE4__SIM_DEVICE    32'h00000052
`define CMACE4__SIM_DEVICE_SZ 152

`define CMACE4__TEST_MODE_PIN_CHAR    32'h00000053
`define CMACE4__TEST_MODE_PIN_CHAR_SZ 40

`endif  // B_CMACE4_DEFINES_VH