// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IBUFDS_IBUFDISABLE_INT_DEFINES_VH
`else
`define B_IBUFDS_IBUFDISABLE_INT_DEFINES_VH

// Look-up table parameters
//

`define IBUFDS_IBUFDISABLE_INT_ADDR_N  5
`define IBUFDS_IBUFDISABLE_INT_ADDR_SZ 32
`define IBUFDS_IBUFDISABLE_INT_DATA_SZ 56

// Attribute addresses
//

`define IBUFDS_IBUFDISABLE_INT__DIFF_TERM    32'h00000000
`define IBUFDS_IBUFDISABLE_INT__DIFF_TERM_SZ 40

`define IBUFDS_IBUFDISABLE_INT__DQS_BIAS    32'h00000001
`define IBUFDS_IBUFDISABLE_INT__DQS_BIAS_SZ 40

`define IBUFDS_IBUFDISABLE_INT__IBUF_LOW_PWR    32'h00000002
`define IBUFDS_IBUFDISABLE_INT__IBUF_LOW_PWR_SZ 40

`define IBUFDS_IBUFDISABLE_INT__IOSTANDARD    32'h00000003
`define IBUFDS_IBUFDISABLE_INT__IOSTANDARD_SZ 56

`define IBUFDS_IBUFDISABLE_INT__USE_IBUFDISABLE    32'h00000004
`define IBUFDS_IBUFDISABLE_INT__USE_IBUFDISABLE_SZ 40

`endif  // B_IBUFDS_IBUFDISABLE_INT_DEFINES_VH