LIBRARY ieee ;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--library work;

entity tb_lane_ctrl_word_insert is
end entity;

architecture tb of tb_lane_ctrl_word_insert is


component lane_ctrl_word_insert is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP

      -- From DATA-LINK/TOP
      RD_DATA_FROM_DL                  : out std_logic;                       --! Read command to receive data from Data-link layer
      CAPABILITY_FROM_DL               : in  std_logic_vector(07 downto 00);  --! Capability field from DATA-LINK layer
      DATA_TX_FROM_DL                  : in  std_logic_vector(31 downto 00);  --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_FROM_DL           : in  std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character from DATA-LINK layer
      NO_DATA_FROM_DL                  : in  std_logic;                       --! Flag to enable the send of IDLE words when no data should be available from Data-Link

      -- From/To skip_insertion
      WAIT_SEND_DATA_FROM_SKIP         : in  std_logic;                       --! Flag to indicates that the skip_insertion send a SKIP control word
      NEW_DATA_TO_SKIP                 : out std_logic;                       --! New data send to skip_insertion
      DATA_TX_TO_SKIP                  : out std_logic_vector(31 downto 00);  --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_TO_SKIP           : out std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character

      -- TX signals command from/to lane_init_fsm
      SEND_INIT1_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT2 control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT3 control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA               : in  std_logic;                       --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS       : in  std_logic;                       --! Flag to send STANDBY control word x32
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  --! Standby reason from MIB
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   : in  std_logic;                       --! Flag to send LOSS_SIGNAL control word x32
      LOST_CAUSE                       : in  std_logic_vector(01 downto 00);  --! Flag to indicate the reason of the LOST_SIGNAL
      STANDBY_SIGNAL_X32               : out std_logic;                       --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32                  : out std_logic                        --! Flag LOST_SIGNAL control word has been send x32
   );
end component;


----------------------------- Stimulus signals
constant periode                       : time := 6.667 ns;

signal RST_N                            : std_logic := '0';
signal CLK                              : std_logic := '0';
-- From DATA-LINK/TOP
signal RD_DATA_FROM_DL                  : std_logic := '0';
signal CAPABILITY_FROM_DL               : std_logic_vector(07 downto 00) := (others => '0');
signal DATA_TX_FROM_DL                  : std_logic_vector(31 downto 00) := (others => '0');
signal VALID_K_CHARAC_FROM_DL           : std_logic_vector(03 downto 00) := (others => '0');
signal NO_DATA_FROM_DL                  : std_logic := '0';
signal WAIT_SEND_DATA_FROM_SKIP         : std_logic := '0';
signal NEW_DATA_TO_SKIP                 : std_logic := '0';
signal DATA_TX_TO_SKIP                  : std_logic_vector(31 downto 00) := (others => '0');
signal VALID_K_CHARAC_TO_SKIP           : std_logic_vector(03 downto 00) := (others => '0');
signal SEND_INIT1_CTRL_WORD             : std_logic := '0';
signal SEND_INIT2_CTRL_WORD             : std_logic := '0';
signal SEND_INIT3_CTRL_WORD             : std_logic := '0';
signal ENABLE_TRANSM_DATA               : std_logic := '0';
signal SEND_32_STANDBY_CTRL_WORDS       : std_logic := '0';
signal STANDBY_REASON                   : std_logic_vector(07 downto 00) := (others => '0');
signal SEND_32_LOSS_SIGNAL_CTRL_WORDS   : std_logic := '0';
signal LOST_CAUSE                       : std_logic_vector(01 downto 00) := (others => '0');
signal STANDBY_SIGNAL_X32               : std_logic := '0';
signal LOST_SIGNAL_X32                  : std_logic := '0';

begin

----------------------------- Instanciation 
DUT : lane_ctrl_word_insert
port map(
   RST_N                            => RST_N,
   CLK                              => CLK,
   RD_DATA_FROM_DL                  => RD_DATA_FROM_DL,
   CAPABILITY_FROM_DL               => CAPABILITY_FROM_DL,
   DATA_TX_FROM_DL                  => DATA_TX_FROM_DL,
   VALID_K_CHARAC_FROM_DL           => VALID_K_CHARAC_FROM_DL,
   NO_DATA_FROM_DL                  => NO_DATA_FROM_DL,
   WAIT_SEND_DATA_FROM_SKIP         => WAIT_SEND_DATA_FROM_SKIP,
   NEW_DATA_TO_SKIP                 => NEW_DATA_TO_SKIP,
   DATA_TX_TO_SKIP                  => DATA_TX_TO_SKIP,
   VALID_K_CHARAC_TO_SKIP           => VALID_K_CHARAC_TO_SKIP,
   SEND_INIT1_CTRL_WORD             => SEND_INIT1_CTRL_WORD,
   SEND_INIT2_CTRL_WORD             => SEND_INIT2_CTRL_WORD,
   SEND_INIT3_CTRL_WORD             => SEND_INIT3_CTRL_WORD,
   ENABLE_TRANSM_DATA               => ENABLE_TRANSM_DATA,
   SEND_32_STANDBY_CTRL_WORDS       => SEND_32_STANDBY_CTRL_WORDS,
   STANDBY_REASON                   => STANDBY_REASON,
   SEND_32_LOSS_SIGNAL_CTRL_WORDS   => SEND_32_LOSS_SIGNAL_CTRL_WORDS,
   LOST_CAUSE                       => LOST_CAUSE,
   STANDBY_SIGNAL_X32               => STANDBY_SIGNAL_X32,
   LOST_SIGNAL_X32                  => LOST_SIGNAL_X32
);


-- generate clock 150 MHz
horloge : process
begin
   CLK   <= not CLK;
   wait for periode/2;
end process;

scenario : process
begin

   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 20 us;
   
   -- Tests of INIT1/2/3
   CAPABILITY_FROM_DL  <= x"FF";
   
   wait until rising_edge(CLK);
   SEND_INIT1_CTRL_WORD <= '1';
   wait for 500 ns;
   wait until rising_edge(CLK);
   SEND_INIT1_CTRL_WORD <= '0';
   SEND_INIT2_CTRL_WORD <= '1';
   wait for 3 us;
   wait until rising_edge(CLK);
   SEND_INIT2_CTRL_WORD <= '0';
   SEND_INIT3_CTRL_WORD <= '1';


   -- Tests active_st no data from DL
   ENABLE_TRANSM_DATA   <= '1';
   NO_DATA_FROM_DL      <= '1';

   --tests active_st data from DL
   --ENABLE_TRANSM_DATA   <= '1';
   --wait until rising_edge(CLK);
   --test_loop : for k in 0 to 50 loop
   --   wait until rising_edge(CLK);
   --   NEW_DATA_FROM_DL    <= '1';
   --   DATA_TX_FROM_DL     <= DATA_TX_FROM_DL+1;
   --   wait until rising_edge(CLK);
   --   NEW_DATA_FROM_DL    <= '0';
   --end loop;

   -- test STANDBY
   SEND_32_STANDBY_CTRL_WORDS <= '1';
   STANDBY_REASON             <= x"FF";
   wait until rising_edge(STANDBY_SIGNAL_X32);
   wait until rising_edge(CLK);
   SEND_32_STANDBY_CTRL_WORDS <= '0';

   -- test LOST_LIGNAL
   --SEND_32_LOSS_SIGNAL_CTRL_WORDS      <= '1';
   --LOST_CAUSE                          <= "11";
   --wait until rising_edge(LOST_SIGNAL_X32);
   --wait until rising_edge(CLK);
   --SEND_32_LOSS_SIGNAL_CTRL_WORDS      <= '0';

   
   
   
   wait;   
end process;

end tb;