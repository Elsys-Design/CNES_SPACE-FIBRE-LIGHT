// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IBUF_IBUFDISABLE_DEFINES_VH
`else
`define B_IBUF_IBUFDISABLE_DEFINES_VH

// Look-up table parameters
//

`define IBUF_IBUFDISABLE_ADDR_N  4
`define IBUF_IBUFDISABLE_ADDR_SZ 32
`define IBUF_IBUFDISABLE_DATA_SZ 144

// Attribute addresses
//

`define IBUF_IBUFDISABLE__IBUF_LOW_PWR    32'h00000000
`define IBUF_IBUFDISABLE__IBUF_LOW_PWR_SZ 40

`define IBUF_IBUFDISABLE__IOSTANDARD    32'h00000001
`define IBUF_IBUFDISABLE__IOSTANDARD_SZ 56

`define IBUF_IBUFDISABLE__SIM_DEVICE    32'h00000002
`define IBUF_IBUFDISABLE__SIM_DEVICE_SZ 144

`define IBUF_IBUFDISABLE__USE_IBUFDISABLE    32'h00000003
`define IBUF_IBUFDISABLE__USE_IBUFDISABLE_SZ 72

`endif  // B_IBUF_IBUFDISABLE_DEFINES_VH