-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/07/2024
--
-- Description : This module implements the lane initialization FSM according to the SpaceFibre standard
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_lane_init_fsm is
  port (
    RST_N                               : in  std_logic;                      --! Global reset signal, Active Low
    CLK                                 : in  std_logic;                      --! Clock generated by the GTY IP
    -- Data-link layer interface
    LANE_RESET_DL                       : in  std_logic;                      --! Lane reset command from the Data-Link layer
    -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
    NO_SIGNAL_PLCWD                     : in  std_logic;                      --! Indicates that no signal is received
    RX_NEW_WORD_PLCWD                   : in  std_logic_vector(1 downto 0);   --! Indicates a new word has been received
    DETECTED_INIT1_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT1 control word has been received
    DETECTED_INIT2_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT2 control word has been received
    DETECTED_INIT3_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT3 control word has been received
    DETECTED_INV_INIT1_PLCWD            : in  std_logic_vector(1 downto 0);   --! Indicates that an inverted INIT1 control word has been received
    DETECTED_INV_INIT2_PLCWD            : in  std_logic_vector(1 downto 0);   --! Indicates that an inverted INIT2 control word has been received
    DETECTED_RXERR_WORD_PLCWD           : in  std_logic_vector(1 downto 0);   --! Indicates that a RXERR control word has been detected
    DETECTED_LOSS_SIGNAL_PLCWD          : in  std_logic_vector(1 downto 0);   --! Flag LOSS_SINGAL control word detected
    DETECTED_STANDBY_PLCWD              : in  std_logic_vector(1 downto 0);   --! Flag STANDBY control word detected
    COMMA_K287_RXED_PLCWD               : in  std_logic_vector(1 downto 0);   --! Flag Comma K28.7 has been received
    SEND_RXERR_PLIF                     : out std_logic_vector(1 downto 0);   --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
    INVERT_RX_BITS_PLIF                 : out std_logic;                      --! Flag to Invert rx bit received
    NO_SIGNAL_DETECTION_ENABLED_PLIF    : out std_logic;                      --! Flag to enable the no signal function
    -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
    STANDBY_SIGNAL_X32_PLCWI            : in  std_logic;                      --! Flag STANDBY control word has been send x32
    LOST_SIGNAL_X32_PLCWI               : in  std_logic;                      --! Flag LOST_SIGNAL control word has been send x32
    SEND_INIT1_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send INIT1 control word following by 64 pseudo-random data words
    SEND_INIT2_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send control word following by 64 pseudo-random data words
    SEND_INIT3_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send control word following by 64 pseudo-random data words
    ENABLE_TRANSM_DATA_PLIF             : out std_logic;                      --! Flag to enable to send data
    SEND_32_STANDBY_CTRL_WORDS_PLIF     : out std_logic;                      --! Flag to send STANDBY control word x32
    SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF : out std_logic;                      --! Flag to send LOSS_SIGNAL control word x32
    LOST_CAUSE_PLIF                     : out std_logic_vector(01 downto 00); --! Flag to indicate the reason of the LOST_SIGNAL
    -- ppl_64_init_hssl (PLIH) interface
    RECEIVER_DISABLED_PLIF              : out std_logic;                      --! Flag to enabled RX function of HSSL IP
    CDR_PLIF                            : out std_logic;                      --! Flag to enabled CDR_PLIF function of HSSL IP
    TRANSMITTER_DISABLED_PLIF           : out std_logic;                      --! Flag to enabled TX fonction of HSSL IP
    -- PARAMETERS and STATUS (MIB interface)
    LANE_START_MIB                      : in  std_logic;                      --! Asserts or de-asserts LaneStart for the lane
    AUTOSTART_MIB                       : in  std_logic;                      --! Asserts or de-asserts AutoStart for the lane
    LANE_RESET_MIB                      : in  std_logic;                      --! Asserts or de-asserts LaneReset for the lane
    LANE_STATE_PLIF                     : out std_logic_vector(03 downto 00); --! Indicates the current state of the Lane Initialization state machine
    RX_ERROR_CNT_PLIF                   : out std_logic_vector(07 downto 00); --! Counter of error detected on the RX link
    RX_ERROR_OVF_PLIF                   : out std_logic                       --! Overflow flag of the RX_ERROR_CNT_PLIF
  );
end ppl_64_lane_init_fsm;

architecture rtl of ppl_64_lane_init_fsm is

---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------

-- Lane Initialisation FSM transition conditions process
   -- Type
type lane_init_fsm_type is (
  CLEAR_LINE_ST,         --! Reset state
  DISABLED_ST,           --! Disabled TX and RX State
  WAIT_ST,               --! Waiting State
  STARTED_ST,            --! Configuration INIT1 State
  INVERT_RX_POLARITY_ST, --! Invert RX polarity in case of detection invert control words
  CONNECTING_ST,         --! Configuration INIT2 State
  CONNECTED_ST,          --! Configuration INIT3 State
  ACTIVE_ST,             --! Transmission Data State
  LOSS_OF_SIGNAL_ST,     --! Error state loss of signal
  PREPARE_STANDBY_ST     --! Error state standby
  );
  -- Signals
signal current_state                : lane_init_fsm_type;                        --! Current state of the Lane Initialisation FSM
signal current_state_r              : lane_init_fsm_type;                        --! Current state registered

-- Lane Initialisation FSM action on state process -------------------------------------------------------------
  -- Constants
constant C_2US_AT_150MHZ            : unsigned(08 downto 00) := "1" & x"2B";     --! 300 x 6.667ns = 2us
  -- Signals
signal clear_line_cnt               : unsigned(08 downto 00);                    --! 2us counter
signal clear_line_done              : std_logic;                                 --! Flag indicates that clear_line_cnt reaches C_2US_AT_150MHZ
signal cdr_i                        : std_logic;                                 --! CDR_PLIF enable command
signal enable_init_cnt              : std_logic;                                 --! enable timeout initialisation counter flag

--RX words counter process -------------------------------------------------------------------------------------
  -- Constants
constant C_MAX_RX_WORDS             : unsigned(13 downto 00) := "11" & x"FFF";   --! 16384 words received
  -- Signals
signal rx_words_cnt                 : unsigned(13 downto 00);                    --! Number of words received counter

-- RX error counter process ------------------------------------------------------------------------------------
  -- Constants
constant C_MAX_RXERR_CTRL_WORDS     : unsigned(07 downto 00) := x"FF";           --! 256 RXERR control words received
  -- Signals
signal rx_error_cnt_i               : unsigned(07 downto 00);                    --! RXERR control words counter
signal rx_error_cnt_ovf_i           : std_logic;                                 --! RXERR overflow flag

-- init_timeout_counter process --------------------------------------------------------------------------------
  -- Constants
constant C_TIME_5000_WORD           : unsigned(12 downto 00) := "0" & x"9C4";    --! 5000 / 2 x 13.334ns = 33.4us
  -- Signals
signal init_timeout_cnt             : unsigned(12 downto 00);                    --! Initialisation timeout counter
signal init_timeout_reaches         : std_logic;                                 --! Flag indicates that init_timeout_cnt reaches C_TIME_5000_WORD

-- Detection 3 consecutive LOST_SIGNAL process -----------------------------------------------------------------
  -- Signals
signal loss_signal_x3_cnt           : unsigned(01 downto 00);                    --! Detection of consecutive LOSS_SIGNAL control words received
signal lost_signal_x3               : std_logic;                                 --! Flag indicates that 3 consecutive LOSS_SIGNAL control word has been received

-- Detection 3 consecutive STANDBY process ---------------------------------------------------------------------
  -- Signals
signal standby_signal_x3_cnt        : unsigned(01 downto 00);                    --! Detection of consecutive STANDBY control words received
signal standby_signal_x3            : std_logic;                                 --! Flag indicates that 3 consecutive STANDBY control word has been received

-- INIT1 detection process -------------------------------------------------------------------------------------
  -- Signals
signal inv_init1_rxed_cnt           : unsigned(01 downto 00);                    --! Detection of the inversed INIT1 counter
signal init1_rxed                   : std_logic;                                 --! Flag indicates that an INIT1 control word has been received
signal init1_rxed_r                 : std_logic;                                 --! init1_rxed registered signal
signal inv_init1_rxed_x3            : std_logic;                                 --! Flag indicates that inv_init1_rxed_cnt reaches 3

-- INIT2 detection process ------------------------------------------------------------------------------------
  -- Signals
signal init2_rxed_cnt               : unsigned(01 downto 00);                    --! Detection of the INIT1 counter
signal inv_init2_rxed_cnt           : unsigned(01 downto 00);                    --! Detection of the inversed INIT1 counter
signal init2_rxed_x3                : std_logic;                                 --! Flag indicates that x3 INIT2 control word has been received
signal inv_init2_rxed_x3            : std_logic;                                 --! Flag indicates that inv_init2_rxed_cnt reaches 3
signal init2_rxed                   : std_logic;                                 --! Flag indicates that INIT2 control word has been received
signal detected_init2_r             : std_logic;                                 --! DETECTED_INIT2_PLCWD registered signal
signal detected_inv_init2_r         : std_logic;                                 --! DETECTED_INV_INIT2_PLCWD registered signal

-- INIT3 detection process ------------------------------------------------------------------------------------
  -- Signals
signal init3_rxed_cnt               : unsigned(01 downto 00);                    --! Detection of the INIT3 counter
signal init3_rxed_x3                : std_logic;                                 --! Flag indicates that x3 INIT3 control word has been received
signal init3_rxed_x3_fw             : std_logic;                                 --! Flag indicates that the third INIT3 control word is received on the first word of the data bus
signal detected_init3_r             : std_logic;                                 --! DETECTED_INIT3_PLCWD registered signal
signal comma_k287_rxed_r            : std_logic;                                 --! COMMA_K287_RXED_PLCWD registered signal

-- Process for detection the reception of 1023 words including the reception of at least on INIT1 or INIT2 without RXERR control words
  -- Constants
constant C_1023_WORDS               : unsigned(09 downto 00) := "11" & x"FF";    --! 1023 words received in STARTED_ST or INVERT_RX_POLARITY_ST
  -- Signals
signal rxed_1023_word_cnt           : unsigned(10 downto 00);                    --! Counter of received words
signal rxed_1023_word               : std_logic;                                 --! Flag indicates that rxed_1023_word_cnt reaches C_1023_WORDS

begin
---------------------------------------------------------
-----                  Assignment                   -----
---------------------------------------------------------
  CDR_PLIF            <= cdr_i;
  RX_ERROR_CNT_PLIF   <= std_logic_vector(rx_error_cnt_i);
  RX_ERROR_OVF_PLIF   <= rx_error_cnt_ovf_i;

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_fsm_lane_init_transition
  --! Lane Initialisation FSM transition conditions process
  ---------------------------------------------------------
  p_fsm_lane_init_transition : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      current_state     <= CLEAR_LINE_ST;
      current_state_r   <= CLEAR_LINE_ST;
    elsif rising_edge(CLK) then
      current_state_r   <= current_state;
      case current_state is
        when CLEAR_LINE_ST         => if clear_line_done = '1' then          -- when 2u counter reaches
                                        current_state  <= DISABLED_ST;
                                      else
                                        current_state  <= CLEAR_LINE_ST;
                                      end if;

        when DISABLED_ST           => if LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then -- When a soft reset appears
                                        current_state  <= CLEAR_LINE_ST;
                                      elsif LANE_START_MIB = '1' or AUTOSTART_MIB = '1' then  -- When a start command is detected
                                        current_state  <= WAIT_ST;
                                      else
                                        current_state  <= DISABLED_ST;
                                      end if;

        when WAIT_ST               => if LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then -- When a soft reset appears
                                        current_state  <= CLEAR_LINE_ST;
                                      elsif LANE_START_MIB = '0' and AUTOSTART_MIB = '0' then -- When a start command is not detected
                                        current_state  <= DISABLED_ST;
                                      elsif LANE_START_MIB = '1' or NO_SIGNAL_PLCWD = '0' then  -- When a start command is detected or signal is received
                                        current_state  <= STARTED_ST;
                                      else
                                        current_state  <= WAIT_ST;
                                      end if;

        when STARTED_ST            => if (lost_signal_x3 = '1' or standby_signal_x3 = '1') or init_timeout_reaches = '1' or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state <= CLEAR_LINE_ST;
                                      elsif inv_init1_rxed_x3 = '1' or inv_init2_rxed_x3 = '1' then
                                        current_state  <= INVERT_RX_POLARITY_ST;
                                      elsif rxed_1023_word = '1' then
                                        current_state  <= CONNECTING_ST;
                                      else
                                        current_state  <= STARTED_ST;
                                      end if;

        when INVERT_RX_POLARITY_ST => if NO_SIGNAL_PLCWD = '1' or init_timeout_reaches = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state  <= CLEAR_LINE_ST;
                                      elsif rxed_1023_word = '1' then
                                        current_state  <= CONNECTING_ST;
                                      else
                                        current_state  <= INVERT_RX_POLARITY_ST;
                                      end if;

        when CONNECTING_ST         => if NO_SIGNAL_PLCWD = '1' or init_timeout_reaches = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state  <= CLEAR_LINE_ST;
                                      elsif init2_rxed_x3 = '1' or init3_rxed_x3 = '1' then
                                        if COMMA_K287_RXED_PLCWD(1) ='1' then
                                          current_state  <= CLEAR_LINE_ST;
                                        else
                                          current_state  <= CONNECTED_ST;
                                        end if;
                                      else
                                        current_state  <= CONNECTING_ST;
                                      end if;

        when CONNECTED_ST          => if NO_SIGNAL_PLCWD = '1' or init_timeout_reaches = '1' or COMMA_K287_RXED_PLCWD(0) ='1' or (COMMA_K287_RXED_PLCWD(0) ='1' and init3_rxed_x3 = '0') or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state  <= CLEAR_LINE_ST;
                                      elsif init3_rxed_x3 = '1' then
                                        if LANE_START_MIB = '0' and AUTOSTART_MIB = '0' and init3_rxed_x3_fw = '1' then
                                          current_state  <= PREPARE_STANDBY_ST;
                                        else
                                          current_state  <= ACTIVE_ST;
                                        end if;
                                      else
                                        current_state  <= CONNECTED_ST;
                                      end if;

        when ACTIVE_ST             => if (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state <= CLEAR_LINE_ST;
                                      elsif LANE_START_MIB = '0' and AUTOSTART_MIB = '0' then
                                        current_state  <= PREPARE_STANDBY_ST;
                                      elsif init1_rxed = '1' or NO_SIGNAL_PLCWD = '1' or rx_error_cnt_ovf_i = '1' then
                                        current_state  <= LOSS_OF_SIGNAL_ST;
                                      else
                                        current_state  <= ACTIVE_ST;
                                      end if;

        when LOSS_OF_SIGNAL_ST     => if LOST_SIGNAL_X32_PLCWI = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state <= CLEAR_LINE_ST;
                                      else
                                        current_state  <= LOSS_OF_SIGNAL_ST;
                                      end if;

        when PREPARE_STANDBY_ST    => if STANDBY_SIGNAL_X32_PLCWI = '1' or (lost_signal_x3 = '1' or standby_signal_x3 = '1') or LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' then
                                        current_state <= CLEAR_LINE_ST;
                                      else
                                        current_state  <= PREPARE_STANDBY_ST;
                                      end if;

        when others                => current_state  <= CLEAR_LINE_ST;
      end case;
    end if;
  end process p_fsm_lane_init_transition;

  ---------------------------------------------------------
  -- Process: p_comb_state
  --! Lane Initialisation FSM action on state process
  ---------------------------------------------------------
   p_comb_state : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         clear_line_cnt                      <= (others => '0');  -- Counter 2us of CLEAR_LINE_ST
         clear_line_done                     <= '0';              -- End condition of CLEAR_LINE_ST
         RECEIVER_DISABLED_PLIF              <= '1';              -- Receiver Disable
         TRANSMITTER_DISABLED_PLIF           <= '1';              -- Transmitter Disabled
         cdr_i                               <= '0';              -- CDR_PLIF Disabled
         SEND_INIT1_CTRL_WORD_PLIF           <= '0';              -- stop send INIT1 control word following by 64 pseudo-random data words
         SEND_INIT2_CTRL_WORD_PLIF           <= '0';              -- stop INIT2 control word following by 64 pseudo-random data words
         SEND_INIT3_CTRL_WORD_PLIF           <= '0';              -- stop INIT3 control word following by 64 pseudo-random data words
         enable_init_cnt                     <= '0';              -- enable timeout initialisation counter
         INVERT_RX_BITS_PLIF                 <= '0';              -- do not invert received bits
         ENABLE_TRANSM_DATA_PLIF             <= '0';              -- enable transimission data and control word from data-link layer
         SEND_32_STANDBY_CTRL_WORDS_PLIF     <= '0';              -- stop 32 STANDBY control words
         SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF <= '0';              -- stop 32 LOSS_SIGNAL control words
         NO_SIGNAL_DETECTION_ENABLED_PLIF    <= '0';              -- No_signal detection function disabled
         LANE_STATE_PLIF                     <= (others => '0');  -- Status of the Lane Init FSM
         LOST_CAUSE_PLIF                     <= (others => '0');  -- LOST_SIGNAL reason

      elsif rising_edge(CLK) then

         if current_state = CLEAR_LINE_ST then

            LANE_STATE_PLIF                     <= x"0"; -- Status of the FSM
            RECEIVER_DISABLED_PLIF              <= '1';  -- Receiver Disable
            TRANSMITTER_DISABLED_PLIF           <= '1';  -- Transmitter Disabled
            cdr_i                               <= '0';  -- CDR_PLIF Disabled
            SEND_INIT1_CTRL_WORD_PLIF           <= '0';  -- Send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '0';  -- Send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '0';  -- Send INIT3 control word following by 64 pseudo-random data words
            enable_init_cnt                     <= '0';  -- disable timeout initialisation counter
            INVERT_RX_BITS_PLIF                 <= '0';  -- do not invert received bits
            ENABLE_TRANSM_DATA_PLIF             <= '0';  -- disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS_PLIF     <= '0';  -- Send 32 STANDBY control words
            SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF <= '0';  -- Send 32 LOSS_SIGNAL control words
            NO_SIGNAL_DETECTION_ENABLED_PLIF    <= '0';  -- No_signal detection function disabled
            LOST_CAUSE_PLIF                     <= "00"; -- Reset

            -- Start counter 2us
            if clear_line_cnt >= C_2US_AT_150MHZ then
               clear_line_done   <= '1';              -- End condition of CLEAR_LINE_ST
            else
               clear_line_cnt    <= clear_line_cnt+1; -- Increment to 1 2us counter
               clear_line_done   <= '0';              -- Reset flag
            end if;

         elsif current_state = DISABLED_ST then

            clear_line_cnt                      <= (others => '0');  -- Reset 2us counter to 0
            LANE_STATE_PLIF                     <= x"1"; -- Status of the FSM
            clear_line_done                     <= '0';  -- Reset 2us flag
            TRANSMITTER_DISABLED_PLIF           <= '1';  -- Transmitter Disabled
            RECEIVER_DISABLED_PLIF              <= '1';  -- Receiver Disabled
            cdr_i                               <= '0';  -- CDR_PLIF Disabled

         elsif current_state = WAIT_ST then

            LANE_STATE_PLIF                     <= x"2";
            RECEIVER_DISABLED_PLIF              <= '0';  -- Receiver Enabled
            TRANSMITTER_DISABLED_PLIF           <= '1';  -- Transmitter Disabled
            cdr_i                               <= '0';  -- CDR_PLIF Disabled
            NO_SIGNAL_DETECTION_ENABLED_PLIF    <= '1';  -- No_signal detection function enabled

         elsif current_state = STARTED_ST then

            LANE_STATE_PLIF                     <= x"3"; -- Status of the FSM
            enable_init_cnt                     <= '1';  -- enable timeout initialisation counter
            TRANSMITTER_DISABLED_PLIF           <= '0';  -- Transmitter Enable
            cdr_i                               <= '1';  -- CDR_PLIF Enable
            SEND_INIT1_CTRL_WORD_PLIF           <= '1';  -- send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = INVERT_RX_POLARITY_ST then

            LANE_STATE_PLIF                     <= x"4"; -- Status of the FSM
            TRANSMITTER_DISABLED_PLIF           <= '0';  -- Transmitter Enable
            cdr_i                               <= '1';  -- CDR_PLIF Enable
            INVERT_RX_BITS_PLIF                 <= '1';  -- invert received bits
            SEND_INIT1_CTRL_WORD_PLIF           <= '1';  -- send INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = CONNECTING_ST then

            LANE_STATE_PLIF                     <= x"5";
            SEND_INIT1_CTRL_WORD_PLIF           <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '1';  -- send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '0';  -- stop INIT3 control word following by 64 pseudo-random data words

         elsif current_state = CONNECTED_ST then

            LANE_STATE_PLIF                     <= x"6"; -- Status of the FSM
            SEND_INIT1_CTRL_WORD_PLIF           <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '0';  -- stop INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '1';  -- send INIT3 control word following by 64 pseudo-random data words

         elsif current_state = ACTIVE_ST then

            LANE_STATE_PLIF                     <= x"7"; -- Status of the FSM
            SEND_INIT1_CTRL_WORD_PLIF           <= '0';  -- stop INIT1 control word following by 64 pseudo-random data words
            SEND_INIT2_CTRL_WORD_PLIF           <= '0';  -- send INIT2 control word following by 64 pseudo-random data words
            SEND_INIT3_CTRL_WORD_PLIF           <= '0';  -- send INIT3 control word following by 64 pseudo-random data words
            enable_init_cnt                     <= '0';  -- disable timeout initialisation counter
            ENABLE_TRANSM_DATA_PLIF             <= '1';  -- enable transimission data and control word from data-link layer

         elsif current_state = PREPARE_STANDBY_ST then

            LANE_STATE_PLIF                     <= x"8"; -- Status of the FSM
            ENABLE_TRANSM_DATA_PLIF             <= '0';  -- Disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS_PLIF     <= '1';  -- send 32 STANDBY control words

         elsif current_state = LOSS_OF_SIGNAL_ST then

            LANE_STATE_PLIF                     <= x"9"; -- Status of the FSM
            ENABLE_TRANSM_DATA_PLIF             <= '0';  -- Disable transimission data and control word from data-link layer
            SEND_32_STANDBY_CTRL_WORDS_PLIF     <= '0';  -- stop 32 STANDBY control words
            SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF <= '1';  -- send 32 LOSS_SIGNAL control words

            -- Reason of the LOST_SIGNAL
            if init1_rxed_r = '1' then
               LOST_CAUSE_PLIF  <= "10";
            elsif rx_error_cnt_ovf_i = '1' then
               LOST_CAUSE_PLIF  <= "01";
            elsif NO_SIGNAL_PLCWD = '1' then
               LOST_CAUSE_PLIF  <= "00";
            end if;

         end if;
      end if;
   end process p_comb_state;

--#######################################################################################--
--------------------------------------- RX processes --------------------------------------
--#######################################################################################--
  ---------------------------------------------------------
  -- Process: p_rx_words_counter
  --! RX words receive counter process
  ---------------------------------------------------------
  p_rx_words_counter : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       rx_words_cnt   <= (others => '0');
    elsif rising_edge(CLK) then
       if RX_NEW_WORD_PLCWD = "11"  and rx_words_cnt < C_MAX_RX_WORDS-1 then    -- when 2 new word are received and lower than 16384 words receive
          rx_words_cnt <= rx_words_cnt + 2;
       elsif (RX_NEW_WORD_PLCWD(0) = '1' or  RX_NEW_WORD_PLCWD(1) = '1') and rx_words_cnt < C_MAX_RX_WORDS then    -- when 1 new word is received and lower than 16384 words receive
          rx_words_cnt <= rx_words_cnt + 1;
       elsif rx_words_cnt >= C_MAX_RX_WORDS then
          rx_words_cnt <= (others => '0');
       end if;
    end if;
  end process p_rx_words_counter;

  ---------------------------------------------------------
  -- Process: p_rxerr_counter
  --!  RX error counter process
  ---------------------------------------------------------
  p_rxerr_counter : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      rx_error_cnt_i          <= (others => '0');
      rx_error_cnt_ovf_i      <= '0';
    elsif rising_edge(CLK) then
      if LANE_RESET_MIB = '1' or LANE_RESET_DL = '1' or current_state = CONNECTED_ST then -- Reset RXERR word counter
         rx_error_cnt_i       <= (others => '0');
         rx_error_cnt_ovf_i   <= '0';
      elsif current_state = ACTIVE_ST then
        -- 16384 words are received and a 2 RXERR control word are detected on the data bus
        if rx_words_cnt >= C_MAX_RX_WORDS and DETECTED_RXERR_WORD_PLCWD = "11" then
          if rx_error_cnt_i = C_MAX_RXERR_CTRL_WORDS then -- Overflow gestion
            rx_error_cnt_ovf_i   <= '1';
            rx_error_cnt_i       <= (others => '1');      -- Lock to the max value 0xFF
          else
            rx_error_cnt_ovf_i   <= '0';
            rx_error_cnt_i       <= rx_error_cnt_i + 1;
          end if;

        -- 16384 words are received and a single RXERR control word is detected on the data bus
        elsif rx_words_cnt >= C_MAX_RX_WORDS and (DETECTED_RXERR_WORD_PLCWD(0) = '1' or DETECTED_RXERR_WORD_PLCWD(1) = '1') then
          rx_error_cnt_i <= rx_error_cnt_i;         -- do not increment RXERR word counter (counter = +1-1)

        -- A single RXERR control word is detected for 16384 words
        elsif rx_words_cnt >= C_MAX_RX_WORDS and rx_error_cnt_i /= x"00" then
          rx_error_cnt_i <= rx_error_cnt_i - 1;

        -- 2 RXERR control word are detected in the data bus
        elsif rx_words_cnt <= C_MAX_RX_WORDS and DETECTED_RXERR_WORD_PLCWD = "11" then
          if (rx_error_cnt_i + 1) = C_MAX_RXERR_CTRL_WORDS then -- Overflow gestion
            rx_error_cnt_ovf_i   <= '1';
            rx_error_cnt_i       <= (others => '1');            -- Lock to the max value 0xFF
          else
            rx_error_cnt_ovf_i   <= '0';
            rx_error_cnt_i       <= rx_error_cnt_i + 2;
          end if;

        -- 1 RXERR control word are detected in the data bus
        elsif rx_words_cnt <= C_MAX_RX_WORDS and (DETECTED_RXERR_WORD_PLCWD(0) = '1' or DETECTED_RXERR_WORD_PLCWD(1) = '1') then
          if rx_error_cnt_i = C_MAX_RXERR_CTRL_WORDS then -- Overflow gestion
            rx_error_cnt_ovf_i   <= '1';
            rx_error_cnt_i       <= (others => '1');      -- Lock to the max value 0xFF
          else
            rx_error_cnt_ovf_i   <= '0';
            rx_error_cnt_i       <= rx_error_cnt_i + 1;
          end if;
        end if;
      end if;
    end if;
  end process p_rxerr_counter;

  ---------------------------------------------------------
  -- Process: p_init_timeout_counter
  --! init_timeout_counter process
  ---------------------------------------------------------
  p_init_timeout_counter : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      init_timeout_cnt     <= (others => '0');
      init_timeout_reaches <= '0';
    elsif rising_edge(CLK) then
      if enable_init_cnt = '1' then                      -- When the initialisation timeout counter is launched (In STARTED_ST)
        if init_timeout_cnt >= C_TIME_5000_WORD then    -- When counter reaches 32us (time to send 5000 words with 5Gbits/s)
          init_timeout_reaches <= '1';
        else
          init_timeout_cnt  <= init_timeout_cnt+1;     -- increment counter
        end if;
      else                                               -- When the initialisation timeout counter is reseted (In ACTIVE_ST and CLEAR_LINE_ST)
        init_timeout_cnt     <= (others => '0');        -- reset counter
        init_timeout_reaches <= '0';                    -- Reset flag timeout
      end if;
    end if;
  end process p_init_timeout_counter;

  ---------------------------------------------------------
  -- Process: p_loss_signal_detection
  --! Detection 3 consecutive LOST_SIGNAL process
  ---------------------------------------------------------
  p_loss_signal_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       lost_signal_x3       <= '0';
       loss_signal_x3_cnt   <= "00";
    elsif rising_edge(CLK) then
      -- if the current_state signal is stable and the FSM is in ACTIVE_ST or LOSS_OF_SIGNAL_ST or PREPARE_STANDBY_ST state
      if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = LOSS_OF_SIGNAL_ST or current_state = PREPARE_STANDBY_ST) then
        if RX_NEW_WORD_PLCWD = "11" and  DETECTED_LOSS_SIGNAL_PLCWD = "11" then -- 2 LOST SIGNAL detected
          if loss_signal_x3_cnt >= "01" then
            lost_signal_x3       <= '1';
            loss_signal_x3_cnt   <= "00";
          else
            lost_signal_x3       <= '0';
            loss_signal_x3_cnt   <= loss_signal_x3_cnt+2;
          end if;
        elsif RX_NEW_WORD_PLCWD(0) = '1' and  DETECTED_LOSS_SIGNAL_PLCWD(0) = '1' then -- 1 LOST SIGNAL detected on the first word
          if loss_signal_x3_cnt >= "10" then
            lost_signal_x3       <= '1';
            loss_signal_x3_cnt   <= "00";
          else
            lost_signal_x3       <= '0';
            loss_signal_x3_cnt   <= loss_signal_x3_cnt+1;
          end if;
        elsif RX_NEW_WORD_PLCWD(1) = '1' and  DETECTED_LOSS_SIGNAL_PLCWD(1) = '1' then -- 1 LOST SIGNAL detected on the second word
          if loss_signal_x3_cnt >= "10" then
            lost_signal_x3       <= '1';
            loss_signal_x3_cnt   <= "00";
          else
            lost_signal_x3       <= '0';
            loss_signal_x3_cnt   <= loss_signal_x3_cnt+1;
          end if;
        else
          lost_signal_x3       <= '0';
          loss_signal_x3_cnt   <= "00";
        end if;
      else
        lost_signal_x3       <= '0';
        loss_signal_x3_cnt   <= "00";
      end if;
    end if;
  end process p_loss_signal_detection;

  ---------------------------------------------------------
  -- Process: p_standby_detection
  --! Detection 3 consecutive STANDBY process
  ---------------------------------------------------------
  p_standby_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      standby_signal_x3       <= '0';
      standby_signal_x3_cnt   <= "00";
    elsif rising_edge(CLK) then
      -- if the current_state signal is stable and the FSM is in ACTIVE_ST or LOSS_OF_SIGNAL_ST or PREPARE_STANDBY_ST state
      if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = LOSS_OF_SIGNAL_ST or current_state = PREPARE_STANDBY_ST) then
        if RX_NEW_WORD_PLCWD = "11" and DETECTED_STANDBY_PLCWD = "11" then -- 2 STANDBY SIGNAL detected
            if standby_signal_x3_cnt >= "01" then
              standby_signal_x3       <= '1';
              standby_signal_x3_cnt   <= "00";
            else
              standby_signal_x3       <= '0';
              standby_signal_x3_cnt   <= standby_signal_x3_cnt+2;
            end if;
        elsif RX_NEW_WORD_PLCWD(0) = '1' and DETECTED_STANDBY_PLCWD(0) = '1' then -- 1 STANDBY SIGNAL detected on the first word
            if standby_signal_x3_cnt >= "10" then
              standby_signal_x3       <= '1';
              standby_signal_x3_cnt   <= "00";
            else
              standby_signal_x3       <= '0';
              standby_signal_x3_cnt   <= standby_signal_x3_cnt+1;
            end if;
        elsif RX_NEW_WORD_PLCWD(1) = '1' and DETECTED_STANDBY_PLCWD(1) = '1' then -- 1 STANDBY SIGNAL detected on the second word
          if standby_signal_x3_cnt >= "10" then
            standby_signal_x3       <= '1';
            standby_signal_x3_cnt   <= "00";
          else
            standby_signal_x3       <= '0';
            standby_signal_x3_cnt   <= standby_signal_x3_cnt+1;
          end if;
        else
          standby_signal_x3          <= '0';
          standby_signal_x3_cnt      <= "00";
        end if;
      else
        standby_signal_x3       <= '0';
        standby_signal_x3_cnt   <= "00";
      end if;
    end if;
  end process p_standby_detection;

  ----------------------------------------
  -- Process: p_inv_init1_detection
  --! INV_INIT1 detection process
  ----------------------------------------
  p_inv_init1_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       inv_init1_rxed_x3    <= '0';
       inv_init1_rxed_cnt   <= "00";
    elsif rising_edge(CLK) then
      -- States for detection of at least one INIT1 is received and no rx error is detected
      if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then
        -- word 1 = INV_INIT1 / word 2 = INV_INIT1
        if DETECTED_INV_INIT1_PLCWD = "11" then
          if inv_init1_rxed_cnt >= "01" then
            inv_init1_rxed_cnt <= "00";
            inv_init1_rxed_x3  <= '1';
          else
            inv_init1_rxed_cnt <= inv_init1_rxed_cnt+2;
            inv_init1_rxed_x3  <= '0';
          end if;

        -- word 1 = INV_INIT1 / word 2 = not RXERR
        elsif DETECTED_INV_INIT1_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if inv_init1_rxed_cnt >= "10" then
            inv_init1_rxed_cnt <= "00";
            inv_init1_rxed_x3  <= '1';
          else
            inv_init1_rxed_cnt <= inv_init1_rxed_cnt+1;
            inv_init1_rxed_x3  <= '0';
          end if;

        -- word 1 = INV_INIT1 / word 2 = RXERR
        elsif DETECTED_INV_INIT1_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if inv_init1_rxed_cnt >= "10" then
            inv_init1_rxed_cnt <= "00";
            inv_init1_rxed_x3  <= '1';
          else
            inv_init1_rxed_cnt <= "00";
            inv_init1_rxed_x3  <= '0';
          end if;

        -- word 1 = not RXERR / word 2 = INV_INIT1
        elsif DETECTED_INV_INIT1_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='0' then
          if inv_init1_rxed_cnt >= "10" then
            inv_init1_rxed_cnt <= "00";
            inv_init1_rxed_x3  <= '1';
          else
            inv_init1_rxed_cnt <= inv_init1_rxed_cnt+1;
            inv_init1_rxed_x3  <= '0';
          end if;

        -- word 1 = RXERR / word 2 = INV_INIT1
        elsif DETECTED_INV_INIT1_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='1' then
          inv_init1_rxed_cnt <= to_unsigned(1,inv_init1_rxed_cnt'length);
          inv_init1_rxed_x3  <= '0';

          -- word 1 = RXERR or word 2 = RXERR
        elsif DETECTED_RXERR_WORD_PLCWD /= "00" then
          inv_init1_rxed_cnt   <= "00";
          inv_init1_rxed_x3    <= '0';
        end if;
      else
        inv_init1_rxed_cnt   <= "00";
        inv_init1_rxed_x3    <= '0';
      end if;
    end if;
  end process p_inv_init1_detection;
  ----------------------------------------
  -- Process: p_init1_detection
  --! INIT1 detection process
  ----------------------------------------
  p_init1_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       init1_rxed           <= '0';
       init1_rxed_r         <= '0';
    elsif rising_edge(CLK) then
      init1_rxed_r <= init1_rxed;
      if current_state = current_state_r and (current_state = ACTIVE_ST or current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then
        -- word 2 = INIT1
        if DETECTED_RXERR_WORD_PLCWD(1) ='1' then
          init1_rxed  <= '0'; -- Transition condition to CONNECTING_ST or LOSS_OF_SIGNAL_ST

        -- word 1 = RXERR and word 2 = INIT1
        elsif DETECTED_RXERR_WORD_PLCWD(0) ='1' and DETECTED_INIT1_PLCWD(1) ='1'then
          init1_rxed <= '1';

        else
          -- word 1 = RXERR
          if DETECTED_RXERR_WORD_PLCWD(0) ='1' then
            init1_rxed <= '0';

          -- word 1 = INIT1 or word 2 = INIT1
          elsif DETECTED_INIT1_PLCWD /= "00" then
            init1_rxed <= '1';
          end if;
        end if;
      else
        init1_rxed  <= '0';
      end if;
    end if;
  end process p_init1_detection;
  ---------------------------------------------------------
  -- Process: p_inv_init2_detection
  --!INV_INIT2 detection process
  ---------------------------------------------------------
  p_inv_init2_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       inv_init2_rxed_x3    <= '0';
       inv_init2_rxed_cnt   <= "00";
    elsif rising_edge(CLK) then
      -- States for detection of at least one INV_INIT2 is received
      if current_state = current_state_r and (current_state = CONNECTING_ST or current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then
        -------------------------
        -- INV_INIT2
        -------------------------
        -- word 1 = INV_INIT2 / word 2 = INV_INIT2
        if DETECTED_INV_INIT2_PLCWD = "11" then
          if inv_init2_rxed_cnt >= "01" then
            inv_init2_rxed_cnt <= "00";
            inv_init2_rxed_x3  <= '1';
          else
            inv_init2_rxed_cnt <= inv_init2_rxed_cnt+2;
            inv_init2_rxed_x3  <= '0';
          end if;

        -- word 1 = INV_INIT2 / word 2 = not RXERR
        elsif DETECTED_INV_INIT2_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if inv_init2_rxed_cnt >= "10" then
            inv_init2_rxed_cnt <= "00";
            inv_init2_rxed_x3  <= '1';
          else
            inv_init2_rxed_cnt <= inv_init2_rxed_cnt+1;
            inv_init2_rxed_x3  <= '0';
          end if;

        -- word 1 = INV_INIT2 / word 2 = RXERR
        elsif DETECTED_INV_INIT2_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if inv_init2_rxed_cnt >= "10" then
            inv_init2_rxed_cnt <= "00";
            inv_init2_rxed_x3  <= '1';
          else
            inv_init2_rxed_cnt <= "00";
            inv_init2_rxed_x3  <= '0';
          end if;

        -- word 1 = not RXERR / word 2 = INV_INIT2
        elsif DETECTED_INV_INIT2_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='0' then
          if inv_init2_rxed_cnt >= "10" then
            inv_init2_rxed_cnt <= "00";
            inv_init2_rxed_x3  <= '1';
          else
            inv_init2_rxed_cnt <= inv_init2_rxed_cnt+1;
            inv_init2_rxed_x3  <= '0';
          end if;

        -- word 1 = RXERR / word 2 = INV_INIT2
        elsif DETECTED_INV_INIT2_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='1' then
          inv_init2_rxed_cnt <= to_unsigned(1,inv_init2_rxed_cnt'length);
          inv_init2_rxed_x3  <= '0';

          -- word 1 = RXERR or word 2 = RXERR
        elsif DETECTED_RXERR_WORD_PLCWD /= "00" then
          inv_init2_rxed_cnt   <= "00";
          inv_init2_rxed_x3    <= '0';
        end if;
      else
        inv_init2_rxed_cnt   <= "00";
        inv_init2_rxed_x3    <= '0';
      end if;
    end if;
  end process p_inv_init2_detection;

  ---------------------------------------------------------
  -- Process: p_init2_detection
  --!INIT2 detection process
  ---------------------------------------------------------
  p_init2_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
        init2_rxed_cnt       <= "00";
        init2_rxed_x3        <= '0';
        init2_rxed           <= '0';
    elsif rising_edge(CLK) then
      -- States for detection of at least one INIT2 is received
      if current_state = current_state_r and (current_state = CONNECTING_ST or current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then
        -------------------------
        -- INIT2
        -------------------------
        -- word 1 = INIT2 / word 2 = INIT2
        if DETECTED_INIT2_PLCWD = "11" then
          init2_rxed <= '1';
          if init2_rxed_cnt >= "01" then
            init2_rxed_cnt <= "00";
            init2_rxed_x3  <= '1';
          else
            init2_rxed_cnt <= init2_rxed_cnt+2;
            init2_rxed_x3  <= '0';
          end if;

        -- word 1 = INIT2 / word 2 = not RXERR
        elsif DETECTED_INIT2_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          init2_rxed <= '1';
          if init2_rxed_cnt >= "10" then
            init2_rxed_cnt <= "00";
            init2_rxed_x3  <= '1';
          else
            init2_rxed_cnt <= init2_rxed_cnt+1;
            init2_rxed_x3  <= '0';
          end if;

        -- word 1 = INIT2 / word 2 = RXERR
        elsif DETECTED_INIT2_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          init2_rxed <= '0';
          if init2_rxed_cnt >= "10" then
            init2_rxed_cnt <= "00";
            init2_rxed_x3  <= '1';
          else
            init2_rxed_cnt <= "00";
            init2_rxed_x3  <= '0';
          end if;

        -- word 1 = not RXERR / word 2 = INIT2
        elsif DETECTED_INIT2_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='0' then
          init2_rxed <= '1';
          if init2_rxed_cnt >= "10" then
            init2_rxed_cnt <= "00";
            init2_rxed_x3  <= '1';
          else
            init2_rxed_cnt <= init2_rxed_cnt+1;
            init2_rxed_x3  <= '0';
          end if;

        -- word 1 = RXERR / word 2 = INIT2
        elsif DETECTED_INIT2_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='1' then
          init2_rxed     <= '0';
          init2_rxed_cnt <= to_unsigned(1,init2_rxed_cnt'length);
          init2_rxed_x3  <= '0';

          -- word 1 = RXERR or word 2 = RXERR
        elsif DETECTED_RXERR_WORD_PLCWD /= "00" then
          init2_rxed_cnt   <= "00";
          init2_rxed_x3    <= '0';
          init2_rxed       <= '0';
        end if;
      else
        init2_rxed       <= '0';
        init2_rxed_cnt   <= "00";
        init2_rxed_x3    <= '0';
      end if;
    end if;
  end process p_init2_detection;

  ---------------------------------------------------------
  -- Process: p_init3_detection
  --!INIT3 detection process
  ---------------------------------------------------------
  p_init3_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
        init3_rxed_cnt    <= "00";
        init3_rxed_x3     <= '0';
        comma_k287_rxed_r <= '0';
        init3_rxed_x3_fw  <= '0';
    elsif rising_edge(CLK) then
      comma_k287_rxed_r <= COMMA_K287_RXED_PLCWD(1);
      init3_rxed_x3_fw  <= '0';
      -- States for detection of at least one INIT3 is received
      if current_state = current_state_r and (current_state = CONNECTING_ST or current_state = CONNECTED_ST) then
        -------------------------
        -- INIT3
        -------------------------
        -- word 1 = INIT3 / word 2 = INIT3
        if DETECTED_INIT3_PLCWD = "11" then
          if init3_rxed_cnt >= "01" then
            init3_rxed_cnt <= "00";
            init3_rxed_x3  <= '1';
          else
            init3_rxed_cnt <= init3_rxed_cnt+2;
            init3_rxed_x3  <= '0';
          end if;

        -- word 1 = INIT3 / word 2 = not RXERR
        elsif DETECTED_INIT3_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if init3_rxed_cnt >= "10" then
            init3_rxed_cnt   <= "00";
            init3_rxed_x3    <= '1';
            init3_rxed_x3_fw <= '1';
          else
            init3_rxed_cnt <= init3_rxed_cnt+1;
            init3_rxed_x3  <= '0';
          end if;

        -- word 1 = INIT3 / word 2 = RXERR
        elsif DETECTED_INIT3_PLCWD(0) = '1' and DETECTED_RXERR_WORD_PLCWD(1) ='0' then
          if init3_rxed_cnt >= "10" then
            init3_rxed_cnt   <= "00";
            init3_rxed_x3    <= '1';
            init3_rxed_x3_fw <= '1';
          else
            init3_rxed_cnt <= "00";
            init3_rxed_x3  <= '0';
          end if;

        -- word 1 = not RXERR / word 2 = INIT3
        elsif DETECTED_INIT3_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='0' then
          if init3_rxed_cnt >= "10" then
            init3_rxed_cnt <= "00";
            init3_rxed_x3  <= '1';
          else
            init3_rxed_cnt <= init3_rxed_cnt+1;
            init3_rxed_x3  <= '0';
          end if;

        -- word 1 = RXERR / word 2 = INIT3
        elsif DETECTED_INIT3_PLCWD(1) = '1' and DETECTED_RXERR_WORD_PLCWD(0) ='1' then
          init3_rxed_cnt <= to_unsigned(1,init3_rxed_cnt'length);
          init3_rxed_x3  <= '0';

          -- word 1 = RXERR or word 2 = RXERR
        elsif DETECTED_RXERR_WORD_PLCWD /= "00" then
          init3_rxed_cnt   <= "00";
          init3_rxed_x3    <= '0';
        end if;
      else
        init3_rxed_cnt   <= "00";
        init3_rxed_x3    <= '0';
      end if;
    end if;
  end process p_init3_detection;

  ---------------------------------------------------------
  -- Process: p_init1_or_init2_detection_without_rx_error
  --!Process for detection the reception of 1023 words including the reception of at least on INIT1 or INIT2 without RXERR control words
  ---------------------------------------------------------
  p_init1_or_init2_detection_without_rx_error : process(CLK,RST_N)
  begin
    if RST_N = '0' then
       rxed_1023_word       <= '0';
       rxed_1023_word_cnt   <= (others => '0');
    elsif rising_edge(CLK) then
      -- if the current_state signal is stable and the FSM is in STARTED_ST or INVERT_ST state
      if current_state = current_state_r and (current_state = STARTED_ST or current_state = INVERT_RX_POLARITY_ST) then
        -- NO RXERR detected
        if DETECTED_RXERR_WORD_PLCWD = "00" then
          -- 2 Words received
          if RX_NEW_WORD_PLCWD = "11" then
            -- 1023 words received without RXERR
            if rxed_1023_word_cnt >= C_1023_WORDS-2 then
              rxed_1023_word_cnt   <= (others => '0');
              if init1_rxed = '1' or init2_rxed = '1'  then
                rxed_1023_word    <= '1';
              else
                rxed_1023_word    <= '0';
              end if;
            else
              rxed_1023_word_cnt   <= rxed_1023_word_cnt+2;
              rxed_1023_word       <= '0';
            end if;
          -- 1 Word received
          elsif RX_NEW_WORD_PLCWD = "01" or RX_NEW_WORD_PLCWD = "01" then
            -- 1023 words received without RXERR
            if rxed_1023_word_cnt >= C_1023_WORDS-1 then
              rxed_1023_word_cnt   <= (others => '0');
              if init1_rxed = '1' or init2_rxed = '1'  then
                rxed_1023_word    <= '1';
              else
                rxed_1023_word    <= '0';
              end if;
            else
              rxed_1023_word_cnt   <= rxed_1023_word_cnt+1;
              rxed_1023_word       <= '0';
            end if;
          end if;

        -- Word 1 = No RXERR and word 2 = RXERR
        elsif DETECTED_RXERR_WORD_PLCWD = "10" then
          if RX_NEW_WORD_PLCWD(0) = '1' then
            -- 1023 words received without RXERR
            if rxed_1023_word_cnt >= C_1023_WORDS-1 then
              rxed_1023_word_cnt   <= (others => '0');
              if init1_rxed = '1' or init2_rxed = '1'  then
                rxed_1023_word    <= '1';
              else
                rxed_1023_word    <= '0';
              end if;
            else
              rxed_1023_word_cnt      <= (others => '0');
              rxed_1023_word          <= '0';
            end if;
          else
            rxed_1023_word_cnt      <= (others => '0');
            rxed_1023_word          <= '0';
          end if;

        -- (word 1 = RXERR and word 2 = No RXERR) or (word 1 = RXERR and word2= RXERR)
        else
          rxed_1023_word_cnt      <= (others => '0');
          rxed_1023_word          <= '0';
        end if;
      else
        rxed_1023_word_cnt   <= (others => '0');
        rxed_1023_word       <= '0';
      end if;
    end if;
  end process p_init1_or_init2_detection_without_rx_error;

  ---------------------------------------------------------
  -- Process: p_send_rx_error_word
  --!RXERR word send to data_link when FSM leave ACTIVE_ST process
  ---------------------------------------------------------
  p_send_rx_error_word : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      SEND_RXERR_PLIF  <= "00";
    elsif rising_edge(CLK) then
      if current_state /= ACTIVE_ST and current_state_r = ACTIVE_ST then   -- when the FSM get out from the ACTIVE_ST
        SEND_RXERR_PLIF  <= "11";                                          -- Send 2 RXERR control words to Data-link layer
      else
        SEND_RXERR_PLIF  <= "00";
      end if;
    end if;
  end process p_send_rx_error_word;
end architecture rtl;
