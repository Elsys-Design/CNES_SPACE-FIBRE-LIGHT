-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 16/07/2025
--
-- Description : This module insert control word in the data flow
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_lane_ctrl_word_insert is
   port (
      RST_N                                : in  std_logic;                                          --! global reset
      CLK                                  : in  std_logic;                                          --! Clock generated by HSSL IP
      -- Data-Link interface
      RD_DATA_EN_PLCWI                     : out std_logic;                                          --! Read command to receive data from Data-link layer
      RD_DATA_VALID_DL                     : in  std_logic;                                          --! Data valid flag from Data-link layer
      CAPABILITY_DL                        : in  std_logic_vector(7 downto 0);                       --! Capability field from DATA-LINK layer
      DATA_TX_DL                           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_DL                    : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character from DATA-LINK layer
      NO_DATA_DL                           : in  std_logic;                                          --! Flag to enable the send of IDLE words when no data should be available from Data-Link
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI                  : in  std_logic;                                          --! Flag to indicates that the skip_insertion send a SKIP control word
      NEW_DATA_PLCWI                       : out std_logic;                                          --! New data send to skip_insertion
      DATA_TX_PLCWI                        : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_PLCWI                 : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character
      -- ppl_64_lane_init_fsm (PLIF) interface
      SEND_INIT1_CTRL_WORD_PLIF            : in  std_logic;                                           --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD_PLIF            : in  std_logic;                                           --! Flag to send INIT2 control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD_PLIF            : in  std_logic;                                           --! Flag to send INIT3 control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA_PLIF              : in  std_logic;                                           --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS_PLIF      : in  std_logic;                                           --! Flag to send STANDBY control word x32
      SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF  : in  std_logic;                                           --! Flag to send LOSS_SIGNAL control word x32
      STANDBY_SIGNAL_X32_PLCWI             : out std_logic;                                          --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32_PLCWI                : out std_logic;                                          --! Flag LOST_SIGNAL control word has been send x32
      -- MIB interface
      STANDBY_REASON_MIB                   : in  std_logic_vector(7 downto 0);                       --! Standby reason from MIB
      LOST_CAUSE_MIB                       : in  std_logic_vector(1 downto 0)                        --! Flag to indicate the reason of the LOST_SIGNAL
   );
end ppl_64_lane_ctrl_word_insert;

architecture rtl of ppl_64_lane_ctrl_word_insert is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------

signal prbs_counter      : unsigned(31 downto 0);
signal send_stdby_cnt    : unsigned(5 downto 0);
signal send_loss_sig_cnt : unsigned(5 downto 0);
signal no_data_dl_r      : std_logic;
begin

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_send_data
-- Description: Align the words so that they are at the beginning of the bus.
---------------------------------------------------------
  p_send_data : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      RD_DATA_EN_PLCWI               <= '0';
      NEW_DATA_PLCWI           <= '0';
      DATA_TX_PLCWI            <= (others => '0');
      VALID_K_CHARAC_PLCWI     <= (others => '0');
      prbs_counter             <= (others => '0');
      send_stdby_cnt           <= (others => '0');
      STANDBY_SIGNAL_X32_PLCWI <= '0';
      send_loss_sig_cnt        <= (others => '0');
      LOST_SIGNAL_X32_PLCWI    <= '0';
      no_data_dl_r             <= '0';
    elsif rising_edge(CLK) then
      no_data_dl_r             <= NO_DATA_DL;
      RD_DATA_EN_PLCWI               <= '0';
      STANDBY_SIGNAL_X32_PLCWI <= '0';
      LOST_SIGNAL_X32_PLCWI    <= '0';
      --------------------------------------
      --      INIT Control Word           --
      --------------------------------------
      if SEND_INIT1_CTRL_WORD_PLIF = '1' or SEND_INIT2_CTRL_WORD_PLIF = '1' or SEND_INIT3_CTRL_WORD_PLIF = '1' then  -- When IP shall sent an INIT control word
        if prbs_counter < C_PRBS_COUNTER_64-1 then  -- PRBS sent
          prbs_counter          <= prbs_counter+2;  -- 2 prbs word
          NEW_DATA_PLCWI        <= '1';
          DATA_TX_PLCWI         <= std_logic_vector(prbs_counter+1) & std_logic_vector(prbs_counter);
          VALID_K_CHARAC_PLCWI  <= x"00";
        elsif prbs_counter = C_PRBS_COUNTER_64-1  then -- INIT insertion
          NEW_DATA_PLCWI        <= '1';
          VALID_K_CHARAC_PLCWI  <= x"10";
          prbs_counter          <= (others => '0');
          if SEND_INIT1_CTRL_WORD_PLIF = '1' then                                -- When INIT1 control word shall be send
            DATA_TX_PLCWI <= C_INIT1_WORD & std_logic_vector(prbs_counter);
          elsif SEND_INIT2_CTRL_WORD_PLIF = '1' then                             -- When INIT2 control word shall be send
            DATA_TX_PLCWI <= C_INIT2_WORD & std_logic_vector(prbs_counter);
          elsif SEND_INIT3_CTRL_WORD_PLIF = '1' then                             -- When INIT3 control word shall be send
            DATA_TX_PLCWI <= CAPABILITY_DL & C_INIT3_WORD & std_logic_vector(prbs_counter);
          end if;
        elsif prbs_counter = C_PRBS_COUNTER_64 then  -- INIT insertion
          NEW_DATA_PLCWI        <= '1';
          VALID_K_CHARAC_PLCWI  <= x"01";
          prbs_counter          <= to_unsigned(1,prbs_counter'length); -- 1 prbs word
          if SEND_INIT1_CTRL_WORD_PLIF = '1' then                           -- When INIT1 control word shall be send
            DATA_TX_PLCWI       <= x"00000000" & C_INIT1_WORD;
          elsif SEND_INIT2_CTRL_WORD_PLIF = '1' then                        -- When INIT2 control word shall be send
            DATA_TX_PLCWI       <= x"00000000" & C_INIT2_WORD;
          elsif SEND_INIT3_CTRL_WORD_PLIF = '1' then                        -- When INIT3 control word shall be send
            DATA_TX_PLCWI       <= x"00000000" & CAPABILITY_DL & C_INIT3_WORD;
          end if;
        end if;
      --------------------------------------
      --   Active state: transmit Data    --
      --------------------------------------
      elsif ENABLE_TRANSM_DATA_PLIF = '1' then -- When the lane_init_fsm is in ACTIVE_ST
        NEW_DATA_PLCWI        <= '1';
        if ((no_data_dl_r = '0' and NO_DATA_DL = '1') or NO_DATA_DL = '0') and WAIT_SEND_DATA_PLSI = '0' then
          RD_DATA_EN_PLCWI          <= '1';
          if RD_DATA_VALID_DL ='1' then
            DATA_TX_PLCWI         <= DATA_TX_DL;
            VALID_K_CHARAC_PLCWI  <= VALID_K_CHARAC_DL;
          else
            DATA_TX_PLCWI         <= C_IDLE_WORD & C_IDLE_WORD;
            VALID_K_CHARAC_PLCWI  <= x"11";
          end if;
        elsif((no_data_dl_r = '0' and NO_DATA_DL = '1') or NO_DATA_DL = '0') and WAIT_SEND_DATA_PLSI = '1' then
          RD_DATA_EN_PLCWI         <= '0';
          if RD_DATA_VALID_DL ='1' then
            DATA_TX_PLCWI         <= DATA_TX_DL;
            VALID_K_CHARAC_PLCWI  <= VALID_K_CHARAC_DL;
          else
            DATA_TX_PLCWI         <= C_IDLE_WORD & C_IDLE_WORD;
            VALID_K_CHARAC_PLCWI  <= x"11";
          end if;
        else -- When no data has been send from DATA-LINK layer
          RD_DATA_EN_PLCWI            <= '1';
          DATA_TX_PLCWI         <= C_IDLE_WORD & C_IDLE_WORD;
          VALID_K_CHARAC_PLCWI  <= x"11";
        end if;
      --------------------------------------
      --      Standby Control Word        --
      --------------------------------------
      elsif SEND_32_STANDBY_CTRL_WORDS_PLIF = '1' then -- When the lane_init_fsm is in PREPARE_STANDBY_ST
        if send_stdby_cnt >= C_X32_SIGNAL then    -- When 32 STANDBY control words has been send
          STANDBY_SIGNAL_X32_PLCWI    <= '1';
          send_stdby_cnt              <= (others => '0');
        elsif send_stdby_cnt < C_X32_SIGNAL then
          STANDBY_SIGNAL_X32_PLCWI    <= '0';
          send_stdby_cnt              <= send_stdby_cnt+2;
          NEW_DATA_PLCWI              <= '1';
          DATA_TX_PLCWI               <= STANDBY_REASON_MIB & C_STANDBY_WORD & STANDBY_REASON_MIB & C_STANDBY_WORD;
          VALID_K_CHARAC_PLCWI        <= x"11";
        end if;
      --------------------------------------
      --    Loss Signal Control Word      --
      --------------------------------------
      elsif SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF = '1' then  -- When the lane_init_fsm is in LOSS_OF_SIGNAL_ST
        if send_loss_sig_cnt >= C_X32_SIGNAL then      -- When 32 LOSS_SIGNAL control words has been send
          LOST_SIGNAL_X32_PLCWI   <= '1';
          send_loss_sig_cnt       <= (others =>'0');
        elsif send_loss_sig_cnt < C_X32_SIGNAL then
          LOST_SIGNAL_X32_PLCWI <= '0';
          send_loss_sig_cnt     <= send_loss_sig_cnt+2;
          NEW_DATA_PLCWI        <= '1';
          DATA_TX_PLCWI         <= "000000" & LOST_CAUSE_MIB & C_LOST_SIG_WORD & "000000" & LOST_CAUSE_MIB & C_LOST_SIG_WORD;
          VALID_K_CHARAC_PLCWI  <= x"11";
        end if;
      else
        NEW_DATA_PLCWI        <= '0';
        DATA_TX_PLCWI         <= (others => '0');
        VALID_K_CHARAC_PLCWI  <= (others => '0');
        prbs_counter          <= (others => '0');
        send_stdby_cnt        <= (others => '0');
        send_loss_sig_cnt     <= (others => '0');
      end if;
    end if;
   end process p_send_data;

end architecture rtl;
