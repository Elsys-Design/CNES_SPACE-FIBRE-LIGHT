----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module describe the Output Buffer & Flow control
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

entity data_out_buff is
  port (
    RST_N                 : in  std_logic;                                    --! global reset
    CLK                   : in  std_logic;                                    --! Clock generated by GTY IP
    -- Link Reset
    LINK_RESET_DLRE       : in std_logic;
    -- AXI-Stream interface
    S_AXIS_ARSTN_NW	      : in std_logic;
		S_AXIS_ACLK_NW	      : in std_logic;
		S_AXIS_TREADY_DL      : out std_logic;
		S_AXIS_TDATA_NW       : in std_logic_vector(C_DATA_LENGTH-1 downto 0);
		S_AXIS_TUSER_NW       : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
		S_AXIS_TLAST_NW       : in std_logic;
		S_AXIS_TVALID_NW      : in std_logic;
    -- DOBUF interface
    VC_READY_DOBUF        : out  std_logic;
    DATA_DOBUF            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
    VALID_K_CHARAC_DOBUF  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
    DATA_VALID_DOBUF      : out  std_logic;
    END_PACKET_DOBUF      : out  std_logic;
    VC_RD_EN_DMAC         : in   std_logic;
    --DDES interface
    M_VAL_DDES            : in std_logic_vector(C_M_SIZE-1 downto 0);
    FCT_FAR_END_DDES      : in std_logic;
    -- PPL interface
    LANE_ACTIVE_ST_PPL    : in std_logic;
    --MIB Interface
    FCT_CC_OVF_DOBUF      : out std_logic;
    CREDIT_VC_DOBUF       : out std_logic;
    VC_CONT_MODE_MIB      : in std_logic
  );
end data_out_buff;

architecture rtl of data_out_buff is
     ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Modules Declaration -----------------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
  component FIFO_DC_AXIS_S is
  	generic (
  		-- Users to add parameters here
      G_DWIDTH                : integer := 36;                                 -- Data bus fifo length
      G_AWIDTH                : integer := 10;                                 -- Address bus fifo length
      G_THRESHOLD_HIGH        : integer := 2**10;                              -- high threshold
      G_THRESHOLD_LOW         : integer := 0;                                  -- low threshold
      -- User parameters ends
      S_AXIS_TDATA_WIDTH	    : integer := 32;                                 -- Data AXIS length
  		S_AXIS_TUSER_WIDTH	    : integer := 4                                   -- User AXIS length
  	);
  	port (
  		-- Users to add ports here
  		aresetn      	        : in std_logic;
  		-- Custom interface master (rd)
  		RD_CLK                  : in  std_logic;                                -- Clock
      RD_DATA                 : out std_logic_vector(G_DWIDTH-1 downto 0);    -- Data read bus
      RD_DATA_EN              : in  std_logic;                                -- Read command
      RD_DATA_VLD             : out std_logic;                                -- Data valid
  		-- STATUS FIFO
      cmd_flush               : in  std_logic;                                -- fifo flush
      STATUS_BUSY_FLUSH       : out std_logic;                                -- fifo is flushing
      STATUS_THRESHOLD_HIGH   : out std_logic;                                -- threshold high reached flag (sur WR_CLK)
      STATUS_THRESHOLD_LOW    : out std_logic;                                -- threshold low reached flag (sur RD_CLK)
      STATUS_FULL             : out std_logic;                                -- full fifo flag (sur WR_CLK)
      STATUS_EMPTY            : out std_logic;                                -- empty fifo flag (sur RD_CLK)
      STATUS_LEVEL_WR         : out std_logic_vector(G_AWIDTH-1 downto 0);    -- Niveau de remplissage de la FIFO (sur WR_CLK)
      STATUS_LEVEL_RD         : out std_logic_vector(G_AWIDTH-1 downto 0) ;   -- Niveau de remplissage de la FIFO (sur RD_CLK)
      -- User ports ends
  		-- Do not modify the ports beyond this line
  		-- Ports of Axi SLAVE Bus Interface S00_AXIS
  		S_AXIS_ACLK             : in std_logic;
  		S_AXIS_TREADY         	: out std_logic;
  		S_AXIS_TDATA          	: in std_logic_vector(C_DATA_LENGTH-1 downto 0);
  		S_AXIS_TUSER          	: in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  		S_AXIS_TLAST          	: in std_logic;
  		S_AXIS_TVALID         	: in std_logic
  	);
  end component;

----------------------------- Declaration signals -----------------------------
type data_in_fsm is (
  IDLE_ST,
  WAIT_END_FLUSH_ST,
  ADD_EEP_ST,
  WAIT_EIP_ST
  );

  signal current_state          : data_in_fsm;
  --Fifo signals
  signal rd_data                : std_logic_vector(C_DATA_LENGTH + C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal rd_data_vld            : std_logic;
  signal status_busy_flush      : std_logic;
  signal status_threshold_high  : std_logic;
  signal status_threshold_low   : std_logic;
  signal status_full            : std_logic;
  signal status_empty           : std_logic;

  signal s_axis_tdata_i         : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal s_axis_tuser_i         : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal s_axis_tlast_i         : std_logic;
  signal s_axis_tvalid_i        : std_logic;
  -- continuous mode
  signal cont_mode_flg          : std_logic;
  signal last_k_char            : std_logic;
  signal cmd_flush              : std_logic;
  --Flow control signals
  signal fct_credit_cnt         : unsigned(C_FCT_CC_SIZE-1 downto 0);
  signal eip_out                : std_logic;
  signal eip_in_req             : std_logic;
  signal eip_in_ack             : std_logic;
  signal eip_in_ack_reg1        : std_logic;
  signal eip_in_ack_reg2        : std_logic;
  signal eip_out_ack            : std_logic;
  signal cnt_eip                : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64
  signal cnt_eip_out            : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64
  signal cnt_eip_in             : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64
  signal cnt_eip_in_reg1        : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64
  signal cnt_eip_in_reg2        : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64
  signal data_out               : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_char_out       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal vc_end_packet          : std_logic;
  signal cnt_word_sent          : unsigned(6-1 downto 0);     -- cnt_word sent, max= 64


begin
---------------------------------------------------------
-----                     Assignation               -----
---------------------------------------------------------

  data_out             <= rd_data(C_DATA_LENGTH-1 downto 0);
  valid_k_char_out     <= rd_data(C_DATA_LENGTH+C_BYTE_BY_WORD_LENGTH-1 downto C_DATA_LENGTH);

  DATA_DOBUF           <= rd_data(C_DATA_LENGTH-1 downto 0);
  VALID_K_CHARAC_DOBUF <= rd_data(C_DATA_LENGTH+C_BYTE_BY_WORD_LENGTH-1 downto C_DATA_LENGTH);
  DATA_VALID_DOBUF     <= rd_data_vld;
  END_PACKET_DOBUF     <= vc_end_packet;

---------------------------------------------------------
-----                     Instanciation             -----
---------------------------------------------------------
  -- FIFO_DC_AXIS_S Instanciation
  ints_fifo_dc_axis_s: FIFO_DC_AXIS_S
  generic map (
    G_DWIDTH              => C_DATA_LENGTH + C_BYTE_BY_WORD_LENGTH,
    G_AWIDTH              => C_OUT_BUF_SIZE,
    G_THRESHOLD_HIGH      => (2**C_OUT_BUF_SIZE)-3,
    G_THRESHOLD_LOW       => 2,
    S_AXIS_TDATA_WIDTH    => C_DATA_LENGTH,
    S_AXIS_TUSER_WIDTH    => C_BYTE_BY_WORD_LENGTH
  )
  port map (
    aresetn               => RST_N,
    RD_CLK                => CLK,
    RD_DATA               => rd_data,
    RD_DATA_EN            => VC_RD_EN_DMAC,
    RD_DATA_VLD           => rd_data_vld,
    cmd_flush             => cmd_flush,
    STATUS_BUSY_FLUSH     => status_busy_flush,
    STATUS_THRESHOLD_HIGH => status_threshold_high,
    STATUS_THRESHOLD_LOW  => status_threshold_low,
    STATUS_FULL           => status_full,
    STATUS_EMPTY          => status_empty,
    STATUS_LEVEL_WR       => open,
    STATUS_LEVEL_RD       => open,
    S_AXIS_ACLK           => S_AXIS_ACLK_NW,
    S_AXIS_TREADY         => S_AXIS_TREADY_DL,
    S_AXIS_TDATA          => s_axis_tdata_i,
    S_AXIS_TUSER          => s_axis_tuser_i,
    S_AXIS_TLAST          => s_axis_tlast_i,
    S_AXIS_TVALID         => s_axis_tvalid_i
  );
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_continuous_mode
-- Description: Manages continuous mode procedure trigger
---------------------------------------------------------
p_continuous_mode: process(CLK, RST_N)
begin
  if RST_N = '0' then
    cont_mode_flg <= '0';
  elsif rising_edge(CLK) then
    cont_mode_flg  <= '0';
    if VC_CONT_MODE_MIB = '1' and (status_threshold_high ='1' or LANE_ACTIVE_ST_PPL ='0') then
        cont_mode_flg  <= '1';
    end if;
  end if;
end process p_continuous_mode;
---------------------------------------------------------
-- Process: p_data_in_fifo
-- Description: Manages the data written into the fifo
---------------------------------------------------------
p_data_in_fifo: process(S_AXIS_ARSTN_NW, S_AXIS_ACLK_NW)
begin
  if S_AXIS_ARSTN_NW = '0' then
    s_axis_tdata_i  <= (others => '0');
    s_axis_tuser_i  <= (others => '0');
    s_axis_tlast_i  <= '0';
    s_axis_tvalid_i <= '0';
    cmd_flush       <= '0';
    current_state   <= IDLE_ST;
  elsif rising_edge(S_AXIS_ACLK_NW) then
    cmd_flush <= '0';
    case current_state is 
      when IDLE_ST =>
                                  if LINK_RESET_DLRE = '1' then
                                    cmd_flush <= '1';
                                    if last_k_char = '1' then
                                      current_state   <= WAIT_END_FLUSH_ST;
                                      s_axis_tdata_i  <= S_AXIS_TDATA_NW;
                                      s_axis_tuser_i  <= S_AXIS_TUSER_NW;
                                      s_axis_tlast_i  <= S_AXIS_TLAST_NW;
                                      s_axis_tvalid_i <= S_AXIS_TVALID_NW;
                                    end if;
                                  elsif cont_mode_flg  = '1' then
                                    cmd_flush <= '1';
                                    if last_k_char = '1' then
                                      current_state   <= ADD_EEP_ST;
                                      s_axis_tdata_i  <= S_AXIS_TDATA_NW;
                                      s_axis_tuser_i  <= S_AXIS_TUSER_NW;
                                      s_axis_tlast_i  <= S_AXIS_TLAST_NW;
                                      s_axis_tvalid_i <= S_AXIS_TVALID_NW;
                                    end if;
                                  else
                                    s_axis_tdata_i  <= S_AXIS_TDATA_NW;
                                    s_axis_tuser_i  <= S_AXIS_TUSER_NW;
                                    s_axis_tlast_i  <= S_AXIS_TLAST_NW;
                                    s_axis_tvalid_i <= S_AXIS_TVALID_NW;
                                  end if;

        when WAIT_END_FLUSH_ST =>
                                  if status_busy_flush = '0' and LINK_RESET_DLRE = '0' then
                                    current_state <= WAIT_EIP_ST;
                                  end if;

        when ADD_EEP_ST =>        if status_busy_flush= '0' and LINK_RESET_DLRE = '0' then
                                    current_state   <= WAIT_EIP_ST;
                                    s_axis_tdata_i  <= C_FILL_SYMB & C_FILL_SYMB & C_FILL_SYMB & C_EEP_SYMB;
                                    s_axis_tuser_i  <= "1111";
                                    s_axis_tlast_i  <= '1';
                                    s_axis_tvalid_i <= '1';
                                  end if;

        when WAIT_EIP_ST =>
                                  if S_AXIS_TUSER_NW(0)='1' and (S_AXIS_TDATA_NW(7 downto 0) = C_EEP_SYMB or S_AXIS_TDATA_NW(7 downto 0) = C_EOP_SYMB) and  S_AXIS_TVALID_NW='1' then
                                    s_axis_tdata_i  <= S_AXIS_TDATA_NW(31 downto 8) & C_FILL_SYMB;
                                    s_axis_tuser_i  <= S_AXIS_TUSER_NW(3 downto 1) & '1';
                                    s_axis_tlast_i  <= '0';
                                    s_axis_tvalid_i <= '1';
                                  elsif S_AXIS_TUSER_NW(1)='1' and (S_AXIS_TDATA_NW(15 downto 8) = C_EEP_SYMB or S_AXIS_TDATA_NW(15 downto 8) = C_EOP_SYMB) and  S_AXIS_TVALID_NW='1' then
                                    s_axis_tdata_i  <= S_AXIS_TDATA_NW(31 downto 16) & C_FILL_SYMB & C_FILL_SYMB;
                                    s_axis_tuser_i  <= S_AXIS_TUSER_NW(3 downto 2) & "11";
                                    s_axis_tlast_i  <= '0';
                                    s_axis_tvalid_i <= '1';
                                  elsif S_AXIS_TUSER_NW(2)='1' and (S_AXIS_TDATA_NW(23 downto 16) = C_EEP_SYMB or S_AXIS_TDATA_NW(23 downto 16) = C_EOP_SYMB) and  S_AXIS_TVALID_NW='1' then
                                    s_axis_tdata_i  <= S_AXIS_TDATA_NW(31 downto 24) & C_FILL_SYMB & C_FILL_SYMB & C_FILL_SYMB;
                                    s_axis_tuser_i  <= S_AXIS_TUSER_NW(3) & "111";
                                    s_axis_tlast_i  <= '0';
                                    s_axis_tvalid_i <= '1';
                                  elsif S_AXIS_TUSER_NW(3)='1' and (S_AXIS_TDATA_NW(31 downto 24) = C_EEP_SYMB or S_AXIS_TDATA_NW(31 downto 24) = C_EOP_SYMB) and  S_AXIS_TVALID_NW='1' then
                                    s_axis_tdata_i  <=  C_FILL_SYMB & C_FILL_SYMB & C_FILL_SYMB & C_FILL_SYMB;
                                    s_axis_tuser_i  <= "1111";
                                    s_axis_tlast_i  <= '0';
                                    s_axis_tvalid_i <= '1';
                                  else
                                    s_axis_tdata_i  <= (others => '0');
                                    s_axis_tuser_i  <= (others => '0');
                                    s_axis_tlast_i  <= '0';
                                    s_axis_tvalid_i <= '0';
                                  end if;
    end case;
  end if;
end process p_data_in_fifo;
---------------------------------------------------------
-- Process: p_last_char_written
-- Description: Analyses if the last character written into
--              the fifo was an EOP, EEP or Fill
---------------------------------------------------------
p_last_char_written: process(S_AXIS_ARSTN_NW, S_AXIS_ACLK_NW)
begin
  if S_AXIS_ARSTN_NW = '0' then
    last_k_char <= '0';
  elsif rising_edge(S_AXIS_ACLK_NW) then
    if S_AXIS_TUSER_NW(C_BYTE_BY_WORD_LENGTH-1)='1' and S_AXIS_TVALID_NW='1' then
      last_k_char <= '1';
    elsif S_AXIS_TVALID_NW='1' then
      last_k_char <= '0';
    end if;
  end if;
end process p_last_char_written;
---------------------------------------------------------
-- Process: p_has_credit
-- Description: Indicates if far end input buffer has credit
---------------------------------------------------------
p_has_credit: process(CLK, RST_N)
begin
  if RST_N = '0' then
    CREDIT_VC_DOBUF <= '0';
  elsif rising_edge(CLK) then
    if fct_credit_cnt > 0 then
      CREDIT_VC_DOBUF <= '1';
    else
      CREDIT_VC_DOBUF <= '0';
    end if;
  end if;
end process p_has_credit;
---------------------------------------------------------
-- Process: p_fct_credit_cnt
-- Description: Manages the FCT credit counter 
---------------------------------------------------------
  p_fct_credit_cnt: process(CLK, RST_N)
  begin
    if RST_N = '0' then
      fct_credit_cnt   <= (others => '0');
      FCT_CC_OVF_DOBUF <= '0';
    elsif rising_edge(CLK) then
      FCT_CC_OVF_DOBUF <= '0';
      if LINK_RESET_DLRE = '1' then
        fct_credit_cnt <= (others => '0');
      else
        if FCT_FAR_END_DDES = '1' and vc_end_packet = '1' then -- FCT received and packet sent
          if C_FCT_CC_MAX > (fct_credit_cnt + (unsigned(M_VAL_DDES)*64)- cnt_word_sent) then -- FCT credit counter will not overflow
            fct_credit_cnt <= fct_credit_cnt + (unsigned(M_VAL_DDES)*64) - cnt_word_sent;
          else
            FCT_CC_OVF_DOBUF <= '1';
            fct_credit_cnt   <= C_FCT_CC_MAX;
          end if;
        elsif vc_end_packet = '1' then -- Packet sent
          if (fct_credit_cnt - cnt_word_sent) > 0 then -- FCT credit counter will not be negative
            fct_credit_cnt <= fct_credit_cnt - cnt_word_sent;
          else
            fct_credit_cnt <= (others => '0');
          end if;
        elsif FCT_FAR_END_DDES = '1' then -- FCT received
          if C_FCT_CC_MAX > fct_credit_cnt + (unsigned(M_VAL_DDES)*64) then -- FCT credit counter will not overflow
           fct_credit_cnt <= fct_credit_cnt + (unsigned(M_VAL_DDES)*64);
          else
            FCT_CC_OVF_DOBUF <= '1';
            fct_credit_cnt   <= C_FCT_CC_MAX;
          end if;
        end if;
      end if;
    end if;
  end process p_fct_credit_cnt;
---------------------------------------------------------
-- Process: p_vc_end_packet
-- Description: EIP output detection
---------------------------------------------------------
p_vc_end_packet: process(CLK, RST_N)
begin
  if RST_N = '0' then
    vc_end_packet <= '0';
  elsif rising_edge(CLK) then
    vc_end_packet <= '0';
    if cnt_word_sent >= 63  and vc_end_packet ='0' then
      vc_end_packet <='1';
    elsif status_threshold_low = '1' and VC_RD_EN_DMAC='1' and vc_end_packet ='0'and cnt_word_sent > 0 then
      vc_end_packet <='1';
    end if;
  end if;
end process p_vc_end_packet;
---------------------------------------------------------
-- Process: p_cnt_word
-- Description: Count the number of word sent
---------------------------------------------------------
p_cnt_word: process(CLK, RST_N)
begin
  if RST_N = '0' then
    cnt_word_sent      <= (others =>'0');
  elsif rising_edge(CLK) then
    if rd_data_vld = '1' and  vc_end_packet='1' then
      cnt_word_sent      <= (others =>'0');
    elsif rd_data_vld = '1' then
      cnt_word_sent <= cnt_word_sent +1;
    elsif cnt_word_sent > 63 then
      cnt_word_sent      <= (others =>'0');
    end if;
  end if;
end process p_cnt_word;
---------------------------------------------------------
-- Process: p_detect_eip_out
-- Description: EIP output detection
---------------------------------------------------------
p_detect_eip_out: process(CLK, RST_N)
begin
  if RST_N = '0' then
    eip_out <= '0';
  elsif rising_edge(CLK) then
    if valid_k_char_out(0)='1' and (data_out(7 downto 0) = C_EEP_SYMB or data_out(7 downto 0) = C_EOP_SYMB) and  VC_RD_EN_DMAC='1' then
      eip_out <= '1';
    elsif valid_k_char_out(1)='1' and (data_out(15 downto 8) = C_EEP_SYMB or data_out(15 downto 8) = C_EOP_SYMB) and  VC_RD_EN_DMAC='1' then
      eip_out <= '1';
    elsif valid_k_char_out(2)='1' and (data_out(23 downto 16) = C_EEP_SYMB or data_out(23 downto 16) = C_EOP_SYMB) and  VC_RD_EN_DMAC='1' then
      eip_out <= '1';
    elsif valid_k_char_out(3)='1' and (data_out(31 downto 24) = C_EEP_SYMB or data_out(31 downto 24) = C_EOP_SYMB) and  VC_RD_EN_DMAC='1' then
      eip_out <= '1';
    else
      eip_out <= '0';
    end if;
  end if;
end process p_detect_eip_out;
---------------------------------------------------------
-- Process: p_eip_cnt
-- Description: Detection of EIP in the buffer
---------------------------------------------------------
p_eip_in: process(S_AXIS_ARSTN_NW, S_AXIS_ACLK_NW)
begin
  if S_AXIS_ARSTN_NW = '0' then
    cnt_eip_in      <= (others =>'0');
    cnt_eip_in_reg1 <= (others =>'0');
    cnt_eip_in_reg2 <= (others =>'0');
    eip_in_req      <= '0';
    eip_in_ack_reg1 <= '0';
    eip_in_ack_reg2 <= '0';
  elsif rising_edge(S_AXIS_ACLK_NW) then
    cnt_eip_in      <= cnt_eip_in;
    cnt_eip_in_reg2 <= cnt_eip_in_reg1;
    eip_in_ack_reg1 <= eip_in_ack;
    eip_in_ack_reg2 <= eip_in_ack_reg1;
    if S_AXIS_TLAST_NW = '1' and eip_in_ack_reg2 ='1' then
      cnt_eip_in <= cnt_eip_in - cnt_eip_in_reg2 + 1;
      eip_in_req <= '0';
    elsif S_AXIS_TLAST_NW = '1' then
      cnt_eip_in <= cnt_eip_in +1;
      eip_in_req <= '1';
    elsif eip_in_ack_reg2 ='1' then
      cnt_eip_in <= cnt_eip_in - cnt_eip_in_reg2;
      eip_in_req <= '0';
    end if;
  end if;
end process p_eip_in;
---------------------------------------------------------
-- Process: p_eip_cnt_out
-- Description: counter of eip in the buffer
---------------------------------------------------------
p_eip_cnt_out: process(CLK, RST_N)
begin
  if RST_N = '0' then
    cnt_eip_out   <= (others =>'0');
  elsif rising_edge(CLK) then
    if eip_out = '1' then
      cnt_eip_out    <= cnt_eip_out + 1;
    elsif eip_out_ack='1' then
      cnt_eip_out   <= (others =>'0');
    end if;
  end if;
end process p_eip_cnt_out;
---------------------------------------------------------
-- Process: p_eip_cnt
-- Description: counter of eip in the buffer
---------------------------------------------------------
p_eip_cnt: process(CLK, RST_N)
begin
  if RST_N = '0' then
    cnt_eip     <= (others =>'0');
    eip_in_ack  <= '0';
    eip_out_ack <= '0';
  elsif rising_edge(CLK) then
    eip_in_ack  <= '0';
    eip_out_ack <= '0';
    if eip_in_req = '1' then
      cnt_eip     <= cnt_eip + cnt_eip_in;
      eip_in_ack  <= '1';
    elsif cnt_eip_out > 0  then
      cnt_eip     <= cnt_eip - cnt_eip_out;
      eip_out_ack <= '1';
    end if;
  end if;
end process p_eip_cnt;
---------------------------------------------------------
-- Process: p_vc_ready
-- Description: Manages the virtual channel ready signal
---------------------------------------------------------
  p_vc_ready: process(CLK, RST_N)
  begin
    if RST_N = '0' then
      VC_READY_DOBUF <= '0';
    elsif rising_edge(CLK) then
      if fct_credit_cnt > 0 and (status_full = '1' or cnt_eip > 0) then
        VC_READY_DOBUF <= '1';
      else
        VC_READY_DOBUF <= '0';
      end if;
    end if;
  end process p_vc_ready;
end architecture rtl;