----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibre_Light Versal target
--
-- Creation date : 03/09/2024
--
-- Description : This module implement the Physical and Lane layer of an IP
-- SpaceFibre Light.
-- The Physical layer is carried by an Xilinx IP
-- The Lane layer is carried by owner's code and an Xilinx IP
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
use phy_plus_lane_lib.pkg_phy_plus_lane.all;

library unisim;
use unisim.vcomponents.all;

library commun;
use commun.all;

entity phy_plus_lane is
   port(
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Main clock
      -- Reset_gen interface 
      LANE_RESET_PPL_OUT               : out std_logic;
      RST_TXCLK_N                      : in  std_logic;                       --! Synchronous reset on clock generated by GTY PLL
      CLK_TX_OUT                       : out std_logic;                       --! Clock generated by manufacturer IP
      RST_TX_DONE                      : out std_logic;                       --! Up when internal rx reset done
      -- CLK GTY signals
      CLK_GTY                          : in std_logic;                        --! Clock for the extended phy layer IP
      -- FROM Data-link layer
      DATA_TX                          : in  std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be send from Data-Link Layer
      LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer
      CAPABILITY_TX                    : in  std_logic_vector(07 downto 00);  --! Capability field send in INIT3 control word
      NEW_DATA_TX                      : in  std_logic;                       --! Flag new data
      VALID_K_CHARAC_TX                : in  std_logic_vector(03 downto 00);  --! 4-bit valid K character flags from Data-link layer
      FIFO_TX_FULL                     : out std_logic;                       --! FiFo TX full flag

      -- TO Data-link layer
      FIFO_RX_RD_EN                    : in  std_logic;                       --! FiFo RX read enable flag
      DATA_RX                          : out std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be received to Data-Link Layer
      FIFO_RX_EMPTY                    : out std_logic;                       --! FiFo RX empty flag
      FIFO_RX_DATA_VALID               : out std_logic;                       --! FiFo RX data valid flag
      VALID_K_CHARAC_RX                : out std_logic_vector(03 downto 00);  --! 4-bit valid K character flags to Data-link layer
      FAR_END_CAPA_DL                  : out std_logic_vector(07 downto 00);  --! Capability field receive in INIT3 control word
      LANE_ACTIVE_DL                   : out std_logic;                       --! Lane Active flag for the DATA Link Layer

      -- FROM/TO Outside
      TX_POS                           : out std_logic;                       --! Positive LVDS serial data send
      TX_NEG                           : out std_logic;                       --! Negative LVDS serial data send
      RX_POS                           : in  std_logic;                       --! Positive LVDS serial data received
      RX_NEG                           : in  std_logic;                       --! Negative LVDS serial data received

      -- PARAMETERS and STATUS
      LANE_START                       : in  std_logic;                       --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                       --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                       --! Asserts or de-asserts LaneReset for the lane
      PARALLEL_LOOPBACK_EN             : in  std_logic;                       --! Enables or disables the parallel loopback for the lane
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  --! In case of error, pauses communication
      NEAR_END_SERIAL_LB_EN            : in  std_logic;                       --! Enables or disables the near-end serial loopback for the lane
      FAR_END_SERIAL_LB_EN             : in  std_logic;                       --! Enables or disables the far-end serial loopback for the lane

      LANE_STATE                       : out std_logic_vector(03 downto 00);  --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic;                       --! Overflow flag of the RX_ERROR_CNT
      LOSS_SIGNAL                      : out std_logic;                       --! Set when no signal is received on RX link
      FAR_END_CAPA                     : out std_logic_vector(07 downto 00);  --! Capabilities field (INT3 flags)
      RX_POLARITY                      : out std_logic                        --! Set when the receiver polarity is inverted
   );
end phy_plus_lane;

architecture rtl of phy_plus_lane is
   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Modules Declaration -----------------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
   component BufG_GT_bd_wrapper is
      port (
        gt_bufgtce_0                      : in  std_logic;
        gt_bufgtcemask_0                  : in  std_logic;
        gt_bufgtclr_0                     : in  std_logic;
        gt_bufgtclrmask_0                 : in  std_logic;
        gt_bufgtdiv_0                     : in  std_logic_vector ( 2 downto 0 );
        outclk_0                          : in  std_logic;
        usrclk_0                          : out std_logic
      );
   end component;

   component FIFO_DC is
      generic (
          G_DWIDTH                : integer := 8;                                 -- Data bus fifo length
          G_AWIDTH                : integer := 8;                                 -- Address bus fifo length
          G_THRESHOLD_HIGH        : integer := 2**8;                              -- high threshold
          G_THRESHOLD_LOW         : integer := 0                                  -- low threshold
      );
      port (
          RST_N                   : in  std_logic;
          -- Writing port
          WR_CLK                  : in  std_logic;                                -- Clock
          WR_DATA                 : in  std_logic_vector(G_DWIDTH-1 downto 0);    -- Data write bus
          WR_DATA_EN              : in  std_logic;                                -- Write command
  
          -- Reading port
          RD_CLK                  : in  std_logic;                                -- Clock
          RD_DATA                 : out std_logic_vector(G_DWIDTH-1 downto 0);    -- Data read bus
          RD_DATA_EN              : in  std_logic;                                -- Read command
          RD_DATA_VLD             : out std_logic;                                -- Data valid
  
          -- Command port
          CMD_FLUSH               : in  std_logic;                                -- fifo flush
          STATUS_BUSY_FLUSH       : out std_logic;                                -- fifo is flushing
  
          -- Status port
          STATUS_THRESHOLD_HIGH   : out std_logic;                                -- threshold high reached flag (sur WR_CLK)
          STATUS_THRESHOLD_LOW    : out std_logic;                                -- threshold low reached flag (sur RD_CLK)
          STATUS_FULL             : out std_logic;                                -- full fifo flag (sur WR_CLK)
          STATUS_EMPTY            : out std_logic;                                -- empty fifo flag (sur RD_CLK)
          STATUS_LEVEL_WR         : out std_logic_vector(G_AWIDTH-1 downto 0);    -- Niveau de remplissage de la FIFO (sur WR_CLK)
          STATUS_LEVEL_RD         : out std_logic_vector(G_AWIDTH-1 downto 0)     -- Niveau de remplissage de la FIFO (sur RD_CLK)
      );
  end component;


   component lane_init_fsm is
      port (
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP
         -- FROM/TO Data-link layer
         LANE_RESET_DL                    : in  std_logic;                       -- Lane reset command from Data-Link Layer.

         -- RX signals
         NO_SIGNAL                        : in  std_logic;                       -- Flag no signal are received
         RX_NEW_WORD                      : in  std_logic;                       -- Flag new word has been received
         DETECTED_INIT1                   : in  std_logic;                       -- Flag INIT1 control word rxed
         DETECTED_INIT2                   : in  std_logic;                       -- Flag INIT2 control word rxed
         DETECTED_INIT3                   : in  std_logic;                       -- Flag INIT3 control word rxed
         DETECTED_INV_INIT1               : in  std_logic;                       -- Flag INV_INIT1 control word rxed
         DETECTED_INV_INIT2               : in  std_logic;                       -- Flag INV_INIT2 control word rxed
         DETECTED_RXERR_WORD              : in  std_logic;                       -- Flag RXERR detected
         DETECTED_LOSS_SIGNAL             : in  std_logic;                       -- Flag LOSS_SINGAL control word detected
         DETECTED_STANDBY                 : in  std_logic;                       -- Flag STANDBY control word detected
         COMMA_K287_RXED                  : in  std_logic;                       -- Flag Comma K28.7 has been received
         RECEIVER_DISABLED                : out std_logic;                       -- flag to enabled RX function of HSSL IP
         CDR                              : out std_logic;                       -- Flag to enabled CDR function of HSSL IP
         SEND_RXERR                       : out std_logic;                       -- Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
         INVERT_RX_BITS                   : out std_logic;                       -- Flag to Invert rx bit received
         NO_SIGNAL_DETECTION_ENABLED      : out std_logic;                       -- Flag to enable the no signal function

         -- TX signals
         STANDBY_SIGNAL_X32               : in  std_logic;                       -- Flag STANDBY control word has been send x32
         LOST_SIGNAL_X32                  : in  std_logic;                       -- Flag LOST_SIGNAL control word has been send x32
         TRANSMITTER_DISABLED             : out std_logic;                       -- flag to enabled TX fonction of HSSL IP
         SEND_INIT1_CTRL_WORD             : out std_logic;                       -- Flag to send INIT1 control word following by 64 pseudo-random data words
         SEND_INIT2_CTRL_WORD             : out std_logic;                       -- Flag to send control word following by 64 pseudo-random data words
         SEND_INIT3_CTRL_WORD             : out std_logic;                       -- Flag to send control word following by 64 pseudo-random data words
         ENABLE_TRANSM_DATA               : out std_logic;                       -- Flag to enable to send data
         SEND_32_STANDBY_CTRL_WORDS       : out std_logic;                       -- Flag to send STANDBY control word x32
         SEND_32_LOSS_SIGNAL_CTRL_WORDS   : out std_logic;                       -- Flag to send LOSS_SIGNAL control word x32
         LOST_CAUSE                       : out std_logic_vector(01 downto 00);  -- Flag to indicate the reason of the LOST_SIGNAL

         -- PARAMETERS and STATUS
         LANE_START                       : in  std_logic;                       -- Asserts or de-asserts LaneStart for the lane
         AUTOSTART                        : in  std_logic;                       -- Asserts or de-asserts AutoStart for the lane
         LANE_RESET                       : in  std_logic;                       -- Asserts or de-asserts LaneReset for the lane
         LANE_STATE                       : out std_logic_vector(03 downto 00);  -- Indicates the current state of the Lane Initialization state machine in a lane
         RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  -- Counter of error detected on the RX link
         RX_ERROR_OVF                     : out std_logic                        -- Overflow flag of the RX_ERROR_CNT
      );
   end component;

   component lane_ctrl_word_insert is
      port (
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP

         -- From DATA-LINK/TOP
         RD_DATA_FROM_DL                  : out std_logic;                       -- Read command to receive data from Data-link layer
         RD_DATA_VALID_FROM_DL            : in  std_logic;                       --! Data valid flag from Data-link layer
         CAPABILITY_FROM_DL               : in  std_logic_vector(07 downto 00);  -- Capability field from DATA-LINK layer
         DATA_TX_FROM_DL                  : in  std_logic_vector(31 downto 00);  -- Data 32-bit receive from DATA_LINK layer
         VALID_K_CHARAC_FROM_DL           : in  std_logic_vector(03 downto 00);  -- Flags indicates which byte is a K character from DATA-LINK layer
         NO_DATA_FROM_DL                  : in  std_logic;                       -- Flag to enable the send of IDLE words when no data should be available from Data-Link
         -- From/To skip_insertion
         WAIT_SEND_DATA_FROM_SKIP         : in  std_logic;                       -- Flag to indicates that the skip_insertion send a SKIP control word
         NEW_DATA_TO_SKIP                 : out std_logic;                       -- New data send to skip_insertion
         DATA_TX_TO_SKIP                  : out std_logic_vector(31 downto 00);  -- Data 32-bit send to manufacturer IP
         VALID_K_CHARAC_TO_SKIP           : out std_logic_vector(03 downto 00);  -- Flags indicates which byte is a K character

         -- TX signals command from/to lane_init_fsm
         SEND_INIT1_CTRL_WORD             : in  std_logic;                       -- Flag to send INIT1 control word following by 64 pseudo-random data words
         SEND_INIT2_CTRL_WORD             : in  std_logic;                       -- Flag to send INIT2 control word following by 64 pseudo-random data words
         SEND_INIT3_CTRL_WORD             : in  std_logic;                       -- Flag to send INIT3 control word following by 64 pseudo-random data words
         ENABLE_TRANSM_DATA               : in  std_logic;                       -- Flag to enable to send data
         SEND_32_STANDBY_CTRL_WORDS       : in  std_logic;                       -- Flag to send STANDBY control word x32
         STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  -- Standby reason from MIB
         SEND_32_LOSS_SIGNAL_CTRL_WORDS   : in  std_logic;                       -- Flag to send LOSS_SIGNAL control word x32
         LOST_CAUSE                       : in  std_logic_vector(01 downto 00);  -- Flag to indicate the reason of the LOST_SIGNAL
         STANDBY_SIGNAL_X32               : out std_logic;                       -- Flag STANDBY control word has been send x32
         LOST_SIGNAL_X32                  : out std_logic                        -- Flag LOST_SIGNAL control word has been send x32
      );
   end component;

   component skip_insertion is
      port (
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP

         -- From/to lane_ctrl_word_insert
         NEW_DATA_FROM_LCWI               : in  std_logic;                       -- New data Flag
         DATA_TX_FROM_LCWI                : in  std_logic_vector(31 downto 00);  -- Data 64-bit receive from DATA_LINK layer
         VALID_K_CHARAC_FROM_LCWI         : in  std_logic_vector(03 downto 00);  -- Flags indicates which byte is a K character from DATA-LINK layer
         WAIT_SEND_DATA                   : out std_logic;                       -- Flag to indicates that the lane_ctrl_word_insert send a SKIP control word

         -- To manufacturer IP
         DATA_TX_TO_IP                    : out std_logic_vector(31 downto 00);  -- Data 64-bit send to manufacturer IP
         VALID_K_CHARAC_TO_IP             : out std_logic_vector(03 downto 00);  -- Flags indicates which byte is a K character

         -- TX signals command from/to lane_init_fsm
         ENABLE_TRANSM_DATA               : in  std_logic                        -- Flag to enable to send data
      );
   end component;

   component parallel_loopback is
      port (
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP
         RST_N                            : in  std_logic;                       -- Global reset
         -- FROM lane_ctrl_word_insert
         DATA_TX_FROM_LCWI                : in  std_logic_vector(31 downto 00);  -- 32-bit Data
         VALID_K_CARAC_FROM_LCWI          : in  std_logic_vector(03 downto 00);  -- 4-bit Valid K character
         DATA_RDY_FROM_LCWI               : in  std_logic;                       -- Data ready flag
         -- FROM rx_sync_fsm
         DATA_TX_FROM_RSF                 : in  std_logic_vector(31 downto 00);  -- 32-bit Data
         VALID_K_CARAC_FROM_RSF           : in  std_logic_vector(03 downto 00);  -- 4-bit Valid K character
         DATA_RDY_FROM_RSF                : in  std_logic;                       -- Data ready flag
         --FROM skip_insertion
         WAIT_SKIP_DATA                   : in  std_logic;                       -- Wait for data to be skip
         --TO lane_ctrl_word_detection
         DATA_TX_TO_LCWD                  : out std_logic_vector(31 downto 00);  -- 32-bit Data
         VALID_K_CARAC_TO_LCWD            : out std_logic_vector(03 downto 00);  -- 4-bit Valid K character
         DATA_RDY_TO_LCWD                 : out std_logic;                       -- Data ready flag
         -- Parameter
         PARALLEL_LOOPBACK_EN             : in  std_logic                        -- Enable or disable the parallel loopback for the lane
      );
   end component;

   component rx_sync_fsm is
      port(
         CLK_SYS                              : in  std_logic;                       --! MAIN CLOCK
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP
         -- FROM Data-link layer
         LANE_RESET_DL                    : in  std_logic;                       -- Lane reset command from Data-Link Layer.
         -- TO lane_ctrl_word_detection
         DATA_RX_TO_LCWD                  : out std_logic_vector(31 downto 00);  -- 32-bit data to lane_ctrl_word_detect
         VALID_K_CARAC_TO_LCWD            : out std_logic_vector(03 downto 00);  -- 4-bit valid K character flags to lane_ctrl_word_detect
         DATA_RDY_TO_LCWD                 : out std_logic;                       -- Data valid flag to lane_ctrl_word_detect
         -- FROM MANUFACTURER IP
         DATA_RX_FROM_IP                  : in  std_logic_vector(31 downto 00);  -- 32-bit data from GTY IP
         VALID_K_CARAC_FROM_IP            : in  std_logic_vector(03 downto 00);  -- 4-bit valid K character flags from GTY IP
         DATA_RDY_FROM_IP                 : in  std_logic;                       -- Data valid flag from GTY IP
         INVALID_CHAR_FROM_IP             : in  std_logic_vector(03 downto 00);  -- Invalid character flags from GTY IP
         DISPARITY_ERR_FROM_IP            : in  std_logic_vector(03 downto 00);  -- Disparity error flags from GTY IP
         RX_WORD_REALIGN_FROM_IP          : in  std_logic;                       -- RX word realign from GTY IP
         COMMA_DET_FROM_IP                : in  std_logic;                       -- Flag indicates that a comma is detected on the word receive
         -- PARAMETERS
         LANE_RESET                       : in  std_logic                        -- Asserts or de-asserts LaneReset for the lane
      );
   end component;

   component lane_ctrl_word_detect is
      port (
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Clock generated by GTY IP

         -- RX control flag signals to from lane_init fsm
         NO_SIGNAL                        : out std_logic;                       -- Flag no signal are received
         RX_NEW_WORD                      : out std_logic;                       -- Flag new word has been received
         DETECTED_INIT1                   : out std_logic;                       -- Flag INIT1 control word rxed
         DETECTED_INIT2                   : out std_logic;                       -- Flag INIT2 control word rxed
         DETECTED_INIT3                   : out std_logic;                       -- Flag INIT3 control word rxed
         DETECTED_INV_INIT1               : out std_logic;                       -- Flag INV_INIT1 control word rxed
         DETECTED_INV_INIT2               : out std_logic;                       -- Flag INV_INIT2 control word rxed
         DETECTED_RXERR_WORD              : out std_logic;                       -- Flag RXERR detected
         DETECTED_LOSS_SIGNAL             : out std_logic;                       -- Flag LOSS_SIGNAL detected
         DETECTED_STANDBY                 : out std_logic;                       -- Flag STANDBY detected
         COMMA_K287_RXED                  : out std_logic;                       -- Flag Comma K28.7 has been received
         CAPABILITY                       : out std_logic_vector(07 downto 00);  -- Capability from INIT3 control word (31 downto 24)
         SEND_RXERR                       : in  std_logic;                       -- Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
         NO_SIGNAL_DETECTION_ENABLED      : in  std_logic;                       -- Flag to enable the no signal function
         ENABLE_TRANSM_DATA               : in  std_logic;                       -- Flag to enable the transmision of data

         -- RX signal from rx_sync_fsm/parallel_loopback
         DATA_RX_FROM_RSF                 : in  std_logic_vector(31 downto 00);  -- 32-bit data from rx_sync_fsm
         VALID_K_CARAC_FROM_RSF           : in  std_logic_vector(03 downto 00);  -- 4-bit valid K character flags from rx_sync_fsm
         DATA_RDY_FROM_RSF                : in  std_logic;                       -- Data valid flag from rx_sync_fsm

         -- RX signals to DATA-LINK
         DATA_RX_TO_DL                    : out std_logic_vector(31 downto 00);  -- 32-bit data to Data-link layer
         VALID_K_CARAC_TO_DL              : out std_logic_vector(03 downto 00);  -- 4-bit valid K character flags to Data-link layer
         DATA_RDY_TO_DL                   : out std_logic                        -- Data valid flag to Data-link layer
      );
   end component;
 component extended_phy_layer_wrapper 
   port (
      INTF0_RX0_ch_rxbufstatus_0 : out STD_LOGIC_VECTOR ( 2 downto 0 );
      INTF0_RX0_ch_rxbyteisaligned_0 : out STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxbyterealign_0 : out STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxcdrhold_0 : in STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxcdrovrden_0 : in STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxcomsasdet_0 : out STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxctrl0_0 : out STD_LOGIC_VECTOR ( 15 downto 0 );
      INTF0_RX0_ch_rxctrl1_0 : out STD_LOGIC_VECTOR ( 15 downto 0 );
      INTF0_RX0_ch_rxctrl2_0 : out STD_LOGIC_VECTOR ( 7 downto 0 );
      INTF0_RX0_ch_rxctrl3_0 : out STD_LOGIC_VECTOR ( 7 downto 0 );
      INTF0_RX0_ch_rxdata_0 : out STD_LOGIC_VECTOR ( 127 downto 0 );
      INTF0_RX0_ch_rxdatavalid_0 : out STD_LOGIC_VECTOR ( 1 downto 0 );
      INTF0_RX0_ch_rxpd_0 : in STD_LOGIC_VECTOR ( 1 downto 0 );
      INTF0_RX0_ch_rxpolarity_0 : in STD_LOGIC_VECTOR ( 0 to 0 );
      INTF0_RX0_ch_rxrate_0 : in STD_LOGIC_VECTOR ( 7 downto 0 );
      INTF0_RX_clr_out_0 : out STD_LOGIC;
      INTF0_RX_clrb_leaf_out_0 : out STD_LOGIC;
      INTF0_TX0_ch_txbufstatus_0 : out STD_LOGIC_VECTOR ( 1 downto 0 );
      INTF0_TX0_ch_txctrl0_0 : in STD_LOGIC_VECTOR ( 15 downto 0 );
      INTF0_TX0_ch_txctrl1_0 : in STD_LOGIC_VECTOR ( 15 downto 0 );
      INTF0_TX0_ch_txctrl2_0 : in STD_LOGIC_VECTOR ( 7 downto 0 );
      INTF0_TX0_ch_txdata : in STD_LOGIC_VECTOR ( 127 downto 0 );
      INTF0_TX0_ch_txpd_0 : in STD_LOGIC_VECTOR ( 1 downto 0 );
      INTF0_TX0_ch_txrate_0 : in STD_LOGIC_VECTOR ( 7 downto 0 );
      INTF0_TX_clr_out_0 : out STD_LOGIC;
      INTF0_TX_clrb_leaf_out_0 : out STD_LOGIC;
      INTF0_rst_all_in_0 : in STD_LOGIC;
      INTF0_rst_rx_datapath_in_0 : in STD_LOGIC;
      INTF0_rst_rx_done_out_0 : out STD_LOGIC;
      INTF0_rst_rx_pll_and_datapath_in_0 : in STD_LOGIC;
      INTF0_rst_tx_datapath_in_0 : in STD_LOGIC;
      INTF0_rst_tx_done_out_0 : out STD_LOGIC;
      INTF0_rst_tx_pll_and_datapath_in_0 : in STD_LOGIC;
      QUAD0_GTREFCLK0_0 : in STD_LOGIC;
      QUAD0_GT_DEBUG_0_gpi : in STD_LOGIC_VECTOR ( 31 downto 0 );
      QUAD0_GT_DEBUG_0_gpo : out STD_LOGIC_VECTOR ( 31 downto 0 );
      QUAD0_RX0_outclk_0 : out STD_LOGIC;
      QUAD0_RX0_usrclk_0 : in STD_LOGIC;
      QUAD0_TX0_outclk_0 : out STD_LOGIC;
      QUAD0_TX0_usrclk_0 : in STD_LOGIC;
      QUAD0_hsclk0_lcplllock_0 : out STD_LOGIC;
      Quad0_CH0_DEBUG_0_ch_loopback : in STD_LOGIC_VECTOR ( 2 downto 0 );
      Quad0_GT_Serial_0_grx_n : in STD_LOGIC_VECTOR ( 3 downto 0 );
      Quad0_GT_Serial_0_grx_p : in STD_LOGIC_VECTOR ( 3 downto 0 );
      Quad0_GT_Serial_0_gtx_n : out STD_LOGIC_VECTOR ( 3 downto 0 );
      Quad0_GT_Serial_0_gtx_p : out STD_LOGIC_VECTOR ( 3 downto 0 );
      gtpowergood_0 : out STD_LOGIC;
      gtwiz_freerun_clk_0 : in STD_LOGIC
    );
 end component;

   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Internal signals declaration --------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
   -- Internal signals from lane_init_fsm
signal transmitter_dis_from_lif                 : std_logic;                        --! Transmitter disable flag from Lane_init_fsm
signal send_init1_ctrl_word_from_lif            : std_logic;                        --! Send INIT1 control word flag from Lane_init_fsm
signal send_init2_ctrl_word_from_lif            : std_logic;                        --! Send INIT2 control word flag from Lane_init_fsm
signal send_init3_ctrl_word_from_lif            : std_logic;                        --! Send INIT3 control word flag from Lane_init_fsm
signal enable_transm_data_from_lif              : std_logic;                        --! Enable transmit data flag from Lane_init_fsm
signal send_32_standby_ctrl_words_from_lif      : std_logic;                        --! Send x32 STANDBY control word flag from Lane_init_fsm
signal send_32_loss_signal_ctrl_word_from_lif   : std_logic;                        --! Send x32 LOSS_SIGNAL control word flag from Lane_init_fsm
signal lost_cause_from_lif                      : std_logic_vector(01 downto 00);   --! LOST cause from Lane_init_fsm
signal lane_state_from_lif                      : std_logic_vector(03 downto 00);   --! Lane state from Lane_init_fsm
signal rx_error_cnt_from_lif                    : std_logic_vector(07 downto 00);   --! RXERR counter from Lane_init_fsm
signal rx_error_ovf_from_lif                    : std_logic;                        --! RXERR counter overflow from Lane_init_fsm
signal receiver_dis_from_lif                    : std_logic;                        --! Receiver disable flag from Lane_init_fsm
signal cdr_from_lif                             : std_logic;                        --! CDR enable from Lane_init_fsm
signal send_rxerr_from_lif                      : std_logic;                        --! Send RXERR control word flag from Lane_init_fsm
signal invert_rx_bits_from_lif                  : std_logic;                        --! RX data invertion flag from Lane_init_fsm
signal no_signal_detection_enabled_from_lif     : std_logic;                        --! No_signal detection enable flag from Lane_init_fsm

   -- Internal signals from FiFos TX
signal data_plus_k_char_from_dl                 : std_logic_vector(35 downto 00);   --! 32-bit Data and 4-bit valid K character from Data_link
signal data_tx_from_fifo                        : std_logic_vector(35 downto 00);   --! 32-bit Data and 4-bit valid K character from TX FiFo
signal fifo_tx_empty                            : std_logic;                        --! TX FiFo empty flag
signal fifo_tx_data_valid                       : std_logic;                        --! TX FiFo data valid flag

   -- Internal signals from lane_ctrl_word_insert
signal rd_data_en_from_lcwi                     : std_logic;                        --! Read data enable flag from Lane_ctrl_word_insert
signal standby_signal_x32_from_lcwi             : std_logic;                        --! x32 STANDBY control words flag (x32 STANDBY has been send) from Lane_ctrl_word_insert
signal lost_signal_x32_from_lcwi                : std_logic;                        --! x32 LOSS_SIGNAL control words flag (x32 LOSS_SIGNAL has been send) from Lane_ctrl_word_insert
signal new_data_from_lcwi                       : std_logic;                        --! New data flag from Lane_ctrl_word_insert
signal data_tx_from_lcwi                        : std_logic_vector(31 downto 00);   --! 32-bit data tx from Lane_ctrl_word_insert
signal valid_k_charac_from_lcwi                 : std_logic_vector(03 downto 00);   --! 4-bit valid K character flags from Lane_ctrl_word_insert

   -- Internal signals from skip_insertion
signal wait_send_data_from_si                   : std_logic;                        --! Wait send data flag from skip_insertion
signal data_tx_from_si                          : std_logic_vector(127 downto 00);  --! 32-bit data from skip_insertion
signal valid_k_charac_from_si                   : std_logic_vector(07 downto 00);   --! 4-bit valid K character flags from skip_insertion

   -- Internal signals from parallel_loopback
signal data_tx_from_plb                         : std_logic_vector(31 downto 00);   --! 32-bit data from parallel_loopback
signal valid_k_charac_from_plb                  : std_logic_vector(03 downto 00);   --! 4-bit valid K character flags from parallel_loopback
signal data_rdy_from_plb                        : std_logic;                        --! Data ready flag from parallel_loopback

   -- Internal signals from rx_sync_fsm
signal data_rx_from_rsf                         : std_logic_vector(31 downto 00);   --! 32-bit data from rx_sync_fsm
signal valid_k_charac_from_rsf                  : std_logic_vector(03 downto 00);   --! 4-bit valid K character flags from rx_sync_fsm
signal data_rdy_from_rsf                        : std_logic;                        --! Data ready flag from rx_sync_fsm

   -- Internal signals from FIFO_RX
signal data_plus_k_char_to_dl                   : std_logic_vector(35 downto 00);   --! 32-bit Data and 4-bit valid K character to Data_link
signal data_plus_k_char_to_fifo_rx              : std_logic_vector(35 downto 00);   --! 32-bit Data and 4-bit valid K character to RX FiFo

   -- Internal signals from lane_ctrl_word_detect
signal no_signal_from_lcwd                      : std_logic;                        --! No_signal flag from lane_ctrl_word_detect
signal rx_new_word_from_lcwd                    : std_logic;                        --! Rx new word receive flag from lane_ctrl_word_detect
signal detected_init1_from_lcwd                 : std_logic;                        --! INIT1 detected flag from lane_ctrl_word_detect
signal detected_init2_from_lcwd                 : std_logic;                        --! INIT2 detected flag from lane_ctrl_word_detect
signal detected_init3_from_lcwd                 : std_logic;                        --! INIT3 detected flag from lane_ctrl_word_detect
signal detected_inv_init1_from_lcwd             : std_logic;                        --! Inversed INIT1 detected flag from lane_ctrl_word_detect
signal detected_inv_init2_from_lcwd             : std_logic;                        --! Inversed INIT2 detected flag from lane_ctrl_word_detect
signal detected_rxerr_word_from_lcwd            : std_logic;                        --! RXERR control word detected flag from lane_ctrl_word_detect
signal detected_lost_signal_from_lcwd           : std_logic;                        --! LOST_SIGNAL control word detected from lane_ctrl_word_detect
signal detected_standby_from_lcwd               : std_logic;                        --! STANDBY control word detected from lane_ctrl_word_detect
signal comma_k287_rxed_from_lcwd                : std_logic;                        --! Comma character K28.7 received flag from lane_ctrl_word_detect
signal data_rx_from_lcwd                        : std_logic_vector(31 downto 00);   --! 32-bit data from lane_ctrl_word_detect
signal valid_k_charac_from_lcwd                 : std_logic_vector(03 downto 00);   --! 4-bit valid K character flags from lane_ctrl_word_detect
signal data_rdy_from_lcwd                       : std_logic;                        --! Data ready flag from lane_ctrl_word_detect
signal far_end_capa_i                           : std_logic_vector(07 downto 00);   --! far_end_capa internal

   -- Internal signals from extended_phy_layer (Manufacturer_IP)
signal QUAD0_TX0_outclk                         : std_logic;                        --! PLL out clock 150MHz generated by GTY IP
signal reset                                    : std_logic;                        --! Reset signal grouping (not RST_N or LANE_RESET or LANE_RESET_DL) in order to reset GTY IP
signal QUAD0_rxp                                : std_logic_vector(03 downto 00);   --! RX positive signal of GTY IP
signal QUAD0_rxn                                : std_logic_vector(03 downto 00);   --! RX negative signal of GTY IP
signal QUAD0_txp                                : std_logic_vector(03 downto 00);   --! TX positive signal of GTY IP
signal QUAD0_txn                                : std_logic_vector(03 downto 00);   --! TX negative signal of GTY IP
signal QUAD0_ch0_loopback                       : std_logic_vector(02 downto 00);   --! Loopback command (Near-end or Far-End loopback) of GTY IP
signal INTF0_RX0_ch_rxcdrhold                   : std_logic_vector(00 downto 00);   --! CRD hold command used in conjunction with INTF0_RX0_ch_rxcdrovrden signal
signal INTF0_RX0_ch_rxcdrovrden                 : std_logic_vector(00 downto 00);   --! CDR Overden command used in conjunction with INTF0_RX0_ch_rxcdrhold signal
signal INTF0_RX0_ch_rxdata                      : std_logic_vector(127 downto 00);  --! 32-bit RX data received and decoded by GTY IP
signal INTF0_RX0_ch_rxdatavalid                 : std_logic_vector(01 downto 00);   --! Data valid flag generated by GTY IP
signal INTF0_RX0_ch_rxbyterealign               : std_logic_vector(00 downto 00);   --! Byte realign flag generated by GTY IP
signal INTF0_RX0_ch_rxctrl0                     : std_logic_vector(15 downto 00);   --! 4-bit valid K character flags generated by GTY IP
signal INTF0_RX0_ch_rxctrl1                     : std_logic_vector(15 downto 00);   --! 4-bit disparity flags generated by GTY IP
signal INTF0_RX0_ch_rxctrl2                     : std_logic_vector(07 downto 00);   --! 4-bit valid comma character flags generated by GTY IP
signal INTF0_RX0_ch_rxctrl3                     : std_logic_vector(07 downto 00);   --! 4-bit not valid charachter flags (in the 8B/10B table) generated by GTY IP
signal QUAD0_hsclk0_lcplllock                   : std_logic;                        --! PLL lock flag generated by the GTY IP
signal INTF0_TX0_ch_txpd                        : std_logic_vector(01 downto 00);   --! Command to disable the transmitter part of GTY IP
signal INTF0_RX0_ch_rxpd                        : std_logic_vector(01 downto 00);   --! Command to disable the receiver part of GTY IP
signal INTF0_rst_tx_done_out_0                  : std_logic;                        --! Up when internal tx reset done
   -- Internal signals from BufG_GT_wrapper
signal clk_tx                                   : std_logic;                        --! Clock generated by the BufG_GT, image of QUAD0_TX0_outclk generated by GTY IP
-- ctrl internal signals
signal ctrl_in_dl               : std_logic_vector(8 downto 0);
signal ctrl_in_dl_sync          : std_logic_vector(8 downto 0);
signal ctrl_out_dl              : std_logic_vector(8 downto 0);
signal ctrl_out_dl_sync         : std_logic_vector(8 downto 0);
signal lane_reset_dl_i          : std_logic;
signal capability_tx_i          : std_logic_vector(7 downto 0);
signal lane_active_dl_i         : std_logic;
signal fifo_in_ctrl_data_valid  : std_logic;
signal fifo_out_ctrl_data_valid : std_logic;
begin

   LANE_RESET_PPL_OUT <= lane_reset_dl_i or LANE_RESET;

   ------------------------------------------------------------------------------
   --! Instance of lane_init_fsm module
   ------------------------------------------------------------------------------
   inst_lane_init_fsm : lane_init_fsm
   port map (
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- FROM/TO Data-link layer
      LANE_RESET_DL                    => lane_reset_dl_i,

      -- RX signals
      NO_SIGNAL                        => no_signal_from_lcwd,
      RX_NEW_WORD                      => rx_new_word_from_lcwd,
      DETECTED_INIT1                   => detected_init1_from_lcwd,
      DETECTED_INIT2                   => detected_init2_from_lcwd,
      DETECTED_INIT3                   => detected_init3_from_lcwd,
      DETECTED_INV_INIT1               => detected_inv_init1_from_lcwd,
      DETECTED_INV_INIT2               => detected_inv_init2_from_lcwd,
      DETECTED_RXERR_WORD              => detected_rxerr_word_from_lcwd,
      DETECTED_LOSS_SIGNAL             => detected_lost_signal_from_lcwd,
      DETECTED_STANDBY                 => detected_standby_from_lcwd,
      COMMA_K287_RXED                  => comma_k287_rxed_from_lcwd,
      RECEIVER_DISABLED                => receiver_dis_from_lif,
      CDR                              => cdr_from_lif,
      SEND_RXERR                       => send_rxerr_from_lif,
      INVERT_RX_BITS                   => invert_rx_bits_from_lif,
      NO_SIGNAL_DETECTION_ENABLED      => no_signal_detection_enabled_from_lif,
      -- TX signals
      STANDBY_SIGNAL_X32               => standby_signal_x32_from_lcwi,
      LOST_SIGNAL_X32                  => lost_signal_x32_from_lcwi,
      TRANSMITTER_DISABLED             => transmitter_dis_from_lif,
      SEND_INIT1_CTRL_WORD             => send_init1_ctrl_word_from_lif,
      SEND_INIT2_CTRL_WORD             => send_init2_ctrl_word_from_lif,
      SEND_INIT3_CTRL_WORD             => send_init3_ctrl_word_from_lif,
      ENABLE_TRANSM_DATA               => enable_transm_data_from_lif,
      SEND_32_STANDBY_CTRL_WORDS       => send_32_standby_ctrl_words_from_lif,
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   => send_32_loss_signal_ctrl_word_from_lif,
      LOST_CAUSE                       => lost_cause_from_lif,
      -- PARAMETERS and STATUS
      LANE_START                       => LANE_START,
      AUTOSTART                        => AUTOSTART,
      LANE_RESET                       => LANE_RESET,
      LANE_STATE                       => lane_state_from_lif,
      RX_ERROR_CNT                     => rx_error_cnt_from_lif,
      RX_ERROR_OVF                     => rx_error_ovf_from_lif
   );
   ------------------------------------------------------------------------------
   -- Instance of TX FIFO_1MB_wrapper module
   ------------------------------------------------------------------------------ 
   ctrl_in_dl      <= LANE_RESET_DL & CAPABILITY_TX;
   lane_reset_dl_i <= '0' when lane_state_from_lif = "0000" else ctrl_in_dl_sync(8) when fifo_in_ctrl_data_valid ='1';
   capability_tx_i <= ctrl_in_dl_sync(7 downto 0) when fifo_in_ctrl_data_valid ='1';
   inst_fifo_in_ctrl : FIFO_DC
   generic map(
        G_DWIDTH                => C_DWIDTH_CTRL_TX,
        G_AWIDTH                => C_AWIDTH_CTRL_TX,
        G_THRESHOLD_HIGH        => 2**C_AWIDTH_CTRL_TX,
        G_THRESHOLD_LOW         => 0
    )
    port map(
        RST_N                   => RST_TXCLK_N,
        -- Writing port
        WR_CLK                  => CLK,
        WR_DATA                 => ctrl_in_dl,
        WR_DATA_EN              => '1',
        -- Reading port
        RD_CLK                  => clk_tx,
        RD_DATA                 => ctrl_in_dl_sync,
        RD_DATA_EN              => '1',
        RD_DATA_VLD             => fifo_in_ctrl_data_valid,
        -- Command port
        CMD_FLUSH               => '0',
        STATUS_BUSY_FLUSH       => open,
        -- Status port
        STATUS_THRESHOLD_HIGH   => open,
        STATUS_THRESHOLD_LOW    => open,
        STATUS_FULL             => open,
        STATUS_EMPTY            => open,
        STATUS_LEVEL_WR         => open,
        STATUS_LEVEL_RD         => open
    );
   ------------------------------------------------------------------------------
   -- Instance of TX FIFO_1MB_wrapper module
   ------------------------------------------------------------------------------ 
   inst_fifo_tx_data : FIFO_DC
   generic map(
        G_DWIDTH                => C_DWIDTH,
        G_AWIDTH                => C_AWIDTH,
        G_THRESHOLD_HIGH        => 2**C_AWIDTH,
        G_THRESHOLD_LOW         => 0
    )
    port map(
        RST_N                   => RST_TXCLK_N,
        -- Writing port
        WR_CLK                  => CLK,
        WR_DATA                 => data_plus_k_char_from_dl,
        WR_DATA_EN              => NEW_DATA_TX,
        -- Reading port
        RD_CLK                  => clk_tx,
        RD_DATA                 => data_tx_from_fifo,
        RD_DATA_EN              => rd_data_en_from_lcwi,
        RD_DATA_VLD             => fifo_tx_data_valid,
        -- Command port
        CMD_FLUSH               => LANE_RESET_DL,
        STATUS_BUSY_FLUSH       => open,
        -- Status port
        STATUS_THRESHOLD_HIGH   => open,
        STATUS_THRESHOLD_LOW    => open,
        STATUS_FULL             => FIFO_TX_FULL,
        STATUS_EMPTY            => fifo_tx_empty,
        STATUS_LEVEL_WR         => open,
        STATUS_LEVEL_RD         => open
    );

   ------------------------------------------------------------------------------
   -- Instance of lane_ctrl_word_insert module
   ------------------------------------------------------------------------------
   inst_lane_ctrl_word_insert : lane_ctrl_word_insert
   port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- From DATA-LINK/TOP
      RD_DATA_FROM_DL                  => rd_data_en_from_lcwi,
      RD_DATA_VALID_FROM_DL            => fifo_tx_data_valid,
      CAPABILITY_FROM_DL               => capability_tx_i,
      DATA_TX_FROM_DL                  => data_tx_from_fifo(31 downto 00),
      VALID_K_CHARAC_FROM_DL           => data_tx_from_fifo(35 downto 32),
      NO_DATA_FROM_DL                  => fifo_tx_empty,
      -- From/To skip_insertion
      WAIT_SEND_DATA_FROM_SKIP         => wait_send_data_from_si,
      NEW_DATA_TO_SKIP                 => new_data_from_lcwi,
      DATA_TX_TO_SKIP                  => data_tx_from_lcwi,
      VALID_K_CHARAC_TO_SKIP           => valid_k_charac_from_lcwi,
      -- TX signals command from/to lane_init_fsm
      SEND_INIT1_CTRL_WORD             => send_init1_ctrl_word_from_lif,
      SEND_INIT2_CTRL_WORD             => send_init2_ctrl_word_from_lif,
      SEND_INIT3_CTRL_WORD             => send_init3_ctrl_word_from_lif,
      ENABLE_TRANSM_DATA               => enable_transm_data_from_lif,
      SEND_32_STANDBY_CTRL_WORDS       => send_32_standby_ctrl_words_from_lif,
      STANDBY_REASON                   => STANDBY_REASON,
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   => send_32_loss_signal_ctrl_word_from_lif,
      LOST_CAUSE                       => lost_cause_from_lif,
      STANDBY_SIGNAL_X32               => standby_signal_x32_from_lcwi,
      LOST_SIGNAL_X32                  => lost_signal_x32_from_lcwi
   );

   ------------------------------------------------------------------------------
   -- Instance of skip_insertion module
   ------------------------------------------------------------------------------
   inst_skip_insertion : skip_insertion
   port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- From/to lane_ctrl_word_insert
      NEW_DATA_FROM_LCWI               => new_data_from_lcwi,
      DATA_TX_FROM_LCWI                => data_tx_from_lcwi,
      VALID_K_CHARAC_FROM_LCWI         => valid_k_charac_from_lcwi,
      WAIT_SEND_DATA                   => wait_send_data_from_si,
      -- To manufacturer IP
      DATA_TX_TO_IP                    => data_tx_from_si(31 downto 00),
      VALID_K_CHARAC_TO_IP             => valid_k_charac_from_si(03 downto 00),
      -- TX signals command from/to lane_init_fsm
      ENABLE_TRANSM_DATA               => enable_transm_data_from_lif
   );

   ------------------------------------------------------------------------------
   -- Instance of parallel_loopback module
   ------------------------------------------------------------------------------
   inst_parallel_loopback : parallel_loopback
   port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- FROM lane_ctrl_word_insert
      DATA_TX_FROM_LCWI                => data_tx_from_lcwi,
      VALID_K_CARAC_FROM_LCWI          => valid_k_charac_from_lcwi,
      DATA_RDY_FROM_LCWI               => new_data_from_lcwi,
      -- FROM rx_sync_fsm
      DATA_TX_FROM_RSF                 => data_rx_from_rsf,
      VALID_K_CARAC_FROM_RSF           => valid_k_charac_from_rsf,
      DATA_RDY_FROM_RSF                => data_rdy_from_rsf,
      -- FROM skip_insertion
      WAIT_SKIP_DATA                   => wait_send_data_from_si,
      --TO lane_ctrl_word_detection
      DATA_TX_TO_LCWD                  => data_tx_from_plb,
      VALID_K_CARAC_TO_LCWD            => valid_k_charac_from_plb,
      DATA_RDY_TO_LCWD                 => data_rdy_from_plb,
      -- Parameter
      PARALLEL_LOOPBACK_EN             => PARALLEL_LOOPBACK_EN
   );


   ------------------------------------------------------------------------------
   -- Instance of rx_sync_fsm module
   ------------------------------------------------------------------------------
   inst_rx_sync_fsm : rx_sync_fsm
   port map(
      CLK_SYS                          => CLK,
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- FROM Data-link layer
      LANE_RESET_DL                    => lane_reset_dl_i,
      -- TO lane_ctrl_word_detection
      DATA_RX_TO_LCWD                  => data_rx_from_rsf,
      VALID_K_CARAC_TO_LCWD            => valid_k_charac_from_rsf,
      DATA_RDY_TO_LCWD                 => data_rdy_from_rsf,
      -- FROM MANUFACTURER IP
      DATA_RX_FROM_IP                  => INTF0_RX0_ch_rxdata(31 downto 00),
      VALID_K_CARAC_FROM_IP            => INTF0_RX0_ch_rxctrl0(03 downto 00),
      DATA_RDY_FROM_IP                 => INTF0_RX0_ch_rxdatavalid(0),
      INVALID_CHAR_FROM_IP             => INTF0_RX0_ch_rxctrl3(03 downto 00),
      DISPARITY_ERR_FROM_IP            => INTF0_RX0_ch_rxctrl1(03 downto 00),
      RX_WORD_REALIGN_FROM_IP          => INTF0_RX0_ch_rxbyterealign(0),
      COMMA_DET_FROM_IP                => INTF0_RX0_ch_rxctrl2(0),
      -- PARAMETERS
      LANE_RESET                       => LANE_RESET
   );

   ------------------------------------------------------------------------------
   -- Instance of lane_ctrl_word_detect module
   ------------------------------------------------------------------------------
   inst_lane_ctrl_word_detect : lane_ctrl_word_detect
   port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- RX control flag signals to from lane_init fsm
      NO_SIGNAL                        => no_signal_from_lcwd,
      RX_NEW_WORD                      => rx_new_word_from_lcwd,
      DETECTED_INIT1                   => detected_init1_from_lcwd,
      DETECTED_INIT2                   => detected_init2_from_lcwd,
      DETECTED_INIT3                   => detected_init3_from_lcwd,
      DETECTED_INV_INIT1               => detected_inv_init1_from_lcwd,
      DETECTED_INV_INIT2               => detected_inv_init2_from_lcwd,
      DETECTED_RXERR_WORD              => detected_rxerr_word_from_lcwd,
      DETECTED_LOSS_SIGNAL             => detected_lost_signal_from_lcwd,
      DETECTED_STANDBY                 => detected_standby_from_lcwd,
      COMMA_K287_RXED                  => comma_k287_rxed_from_lcwd,
      CAPABILITY                       => far_end_capa_i,
      SEND_RXERR                       => send_rxerr_from_lif,
      NO_SIGNAL_DETECTION_ENABLED      => no_signal_detection_enabled_from_lif,
      ENABLE_TRANSM_DATA               => enable_transm_data_from_lif,
      -- RX signal from rx_sync_fsm/parallel_loopback
      DATA_RX_FROM_RSF                 => data_tx_from_plb,
      VALID_K_CARAC_FROM_RSF           => valid_k_charac_from_plb,
      DATA_RDY_FROM_RSF                => data_rdy_from_plb,
      -- RX signals to DATA-LINK
      DATA_RX_TO_DL                    => data_rx_from_lcwd,
      VALID_K_CARAC_TO_DL              => valid_k_charac_from_lcwd,
      DATA_RDY_TO_DL                   => data_rdy_from_lcwd

   );

   ------------------------------------------------------------------------------
   -- Instance of RX FIFO_1MB_wrapper module
   ------------------------------------------------------------------------------
   data_plus_k_char_to_fifo_rx   <= valid_k_charac_from_lcwd & data_rx_from_lcwd;   -- regroup data and valid K char on 36-bit vector

   inst_fifo_rx_data : FIFO_DC
      generic map(
           G_DWIDTH                => C_DWIDTH,
           G_AWIDTH                => C_AWIDTH,
           G_THRESHOLD_HIGH        => 2**C_AWIDTH,
           G_THRESHOLD_LOW         => 0
       )
       port map(
           RST_N                   => RST_N,
           -- Writing port
           WR_CLK                  => clk_tx,
           WR_DATA                 => data_plus_k_char_to_fifo_rx,
           WR_DATA_EN              => data_rdy_from_lcwd,
           -- Reading port
           RD_CLK                  => CLK,
           RD_DATA                 => data_plus_k_char_to_dl,
           RD_DATA_EN              => FIFO_RX_RD_EN,
           RD_DATA_VLD             => FIFO_RX_DATA_VALID,
           -- Command port
           CMD_FLUSH               => LANE_RESET_DL,
           STATUS_BUSY_FLUSH       => open,
           -- Status port
           STATUS_THRESHOLD_HIGH   => open,
           STATUS_THRESHOLD_LOW    => open,
           STATUS_FULL             => open,
           STATUS_EMPTY            => FIFO_RX_EMPTY,
           STATUS_LEVEL_WR         => open,
           STATUS_LEVEL_RD         => open
       );
   ------------------------------------------------------------------------------
   -- Instance of TX FIFO_1MB_wrapper module
   ------------------------------------------------------------------------------ 
   ctrl_out_dl     <= lane_active_dl_i & far_end_capa_i;
   LANE_ACTIVE_DL  <= ctrl_out_dl_sync(8)          when fifo_out_ctrl_data_valid ='1';
   FAR_END_CAPA_DL <= ctrl_out_dl_sync(7 downto 0) when fifo_out_ctrl_data_valid ='1';
   inst_fifo_out_ctrl : FIFO_DC
   generic map(
        G_DWIDTH                => C_DWIDTH_CTRL_RX,
        G_AWIDTH                => C_AWIDTH_CTRL_RX,
        G_THRESHOLD_HIGH        => 2**C_AWIDTH_CTRL_RX,
        G_THRESHOLD_LOW         => 0
    )
    port map(
        RST_N                   => RST_N,
        -- Writing port
        WR_CLK                  => clk_tx,
        WR_DATA                 => ctrl_out_dl,
        WR_DATA_EN              => '1',
        -- Reading port
        RD_CLK                  => CLK,
        RD_DATA                 => ctrl_out_dl_sync,
        RD_DATA_EN              => '1',
        RD_DATA_VLD             => fifo_out_ctrl_data_valid,
        -- Command port
        CMD_FLUSH               => '0',
        STATUS_BUSY_FLUSH       => open,
        -- Status port
        STATUS_THRESHOLD_HIGH   => open,
        STATUS_THRESHOLD_LOW    => open,
        STATUS_FULL             => open,
        STATUS_EMPTY            => open,
        STATUS_LEVEL_WR         => open,
        STATUS_LEVEL_RD         => open
    );
   ------------------------------------------------------------------------------
   -- Instance of TX BufG_GT_wrapper module for TX clock
   ------------------------------------------------------------------------------
      inst_bufg_gt_tx_clock : BufG_GT_bd_wrapper
         port map(
           gt_bufgtce_0                   => '1',
           gt_bufgtcemask_0               => '0',
           gt_bufgtclr_0                  => '0',
           gt_bufgtclrmask_0              => '0',
           gt_bufgtdiv_0                  => "000",
           outclk_0                       => QUAD0_TX0_outclk,
           usrclk_0                       => clk_tx
         );

   reset <= not RST_N or LANE_RESET or lane_reset_dl_i;

   -- Near-End and Far-End loopback drivin function
   QUAD0_ch0_loopback         <= "010"    when NEAR_END_SERIAL_LB_EN = '1' else
                                 "100"    when FAR_END_SERIAL_LB_EN = '1'  else
                                 "000";

   -- Clock Data recovery drivin function
   INTF0_RX0_ch_rxcdrhold     <= "0"      when cdr_from_lif = '1' else "1";
   INTF0_RX0_ch_rxcdrovrden   <= "0"      when cdr_from_lif = '1' else "0";

   -- Disable transmitter and/or receiver drinvin function
   INTF0_TX0_ch_txpd          <= "11"     when transmitter_dis_from_lif = '1' else "00";
   INTF0_RX0_ch_rxpd          <= "11"     when receiver_dis_from_lif = '1' else "00";

   ------------------------------------------------------------------------------
   -- Instance of extended_phy_layer module
   ------------------------------------------------------------------------------
  inst_extended_phy_layer_wrapper : extended_phy_layer_wrapper
   port map(
     INTF0_RX0_ch_rxbufstatus_0           => open,
     INTF0_RX0_ch_rxbyteisaligned_0       => open,
     INTF0_RX0_ch_rxbyterealign_0         => INTF0_RX0_ch_rxbyterealign,
     INTF0_RX0_ch_rxcdrhold_0             => INTF0_RX0_ch_rxcdrhold,
     INTF0_RX0_ch_rxcdrovrden_0           => INTF0_RX0_ch_rxcdrovrden,
     INTF0_RX0_ch_rxcomsasdet_0           => open,
     INTF0_RX0_ch_rxctrl0_0               => INTF0_RX0_ch_rxctrl0,
     INTF0_RX0_ch_rxctrl1_0               => INTF0_RX0_ch_rxctrl1,
     INTF0_RX0_ch_rxctrl2_0               => INTF0_RX0_ch_rxctrl2,
     INTF0_RX0_ch_rxctrl3_0               => INTF0_RX0_ch_rxctrl3,
     INTF0_RX0_ch_rxdata_0                => INTF0_RX0_ch_rxdata,
     INTF0_RX0_ch_rxdatavalid_0           => INTF0_RX0_ch_rxdatavalid,
     INTF0_RX0_ch_rxpd_0                  => INTF0_RX0_ch_rxpd,
     INTF0_RX0_ch_rxpolarity_0(0)         => invert_rx_bits_from_lif,
     INTF0_RX0_ch_rxrate_0                => "00000000",
     INTF0_RX_clr_out_0                   => open,
     INTF0_RX_clrb_leaf_out_0             => open,
     INTF0_TX0_ch_txbufstatus_0           => open,
     INTF0_TX0_ch_txctrl0_0               => "0000000000000000",
     INTF0_TX0_ch_txctrl1_0               => "0000000000000000",
     INTF0_TX0_ch_txctrl2_0               => valid_k_charac_from_si,
     INTF0_TX0_ch_txdata                  => data_tx_from_si,
     INTF0_TX0_ch_txpd_0                  => INTF0_TX0_ch_txpd,
     INTF0_TX0_ch_txrate_0                => "00000000",
     INTF0_TX_clr_out_0                   => open,
     INTF0_TX_clrb_leaf_out_0             => open,
     INTF0_rst_all_in_0                   => reset,
     INTF0_rst_rx_datapath_in_0           => '0',
     INTF0_rst_rx_done_out_0              => open,
     INTF0_rst_rx_pll_and_datapath_in_0   => '0',
     INTF0_rst_tx_datapath_in_0           => '0',
     INTF0_rst_tx_done_out_0              => INTF0_rst_tx_done_out_0,
     INTF0_rst_tx_pll_and_datapath_in_0   => '0',
     QUAD0_GTREFCLK0_0                    => CLK_GTY,
     QUAD0_GT_DEBUG_0_gpi                 => x"00000000",
     QUAD0_GT_DEBUG_0_gpo                 => open,
     QUAD0_RX0_outclk_0                   => open,
     QUAD0_RX0_usrclk_0                   => clk_tx,--QUAD0_TX0_outclk,
     QUAD0_TX0_outclk_0                   => QUAD0_TX0_outclk,
     QUAD0_TX0_usrclk_0                   => clk_tx, --QUAD0_TX0_outclk,
     QUAD0_hsclk0_lcplllock_0             => QUAD0_hsclk0_lcplllock,
     Quad0_CH0_DEBUG_0_ch_loopback        => QUAD0_ch0_loopback,
     Quad0_GT_Serial_0_grx_n              => QUAD0_rxn,
     Quad0_GT_Serial_0_grx_p              => QUAD0_rxp,
     Quad0_GT_Serial_0_gtx_n              => QUAD0_txn,
     Quad0_GT_Serial_0_gtx_p              => QUAD0_txp,
     gtpowergood_0                        => open,
     gtwiz_freerun_clk_0                  => CLK
   );



  -- Inputs/Outputs
CLK_TX_OUT                 <= clk_tx;

data_plus_k_char_from_dl   <= VALID_K_CHARAC_TX & DATA_TX;
DATA_RX                    <= data_plus_k_char_to_dl(31 downto 00);
VALID_K_CHARAC_RX          <= data_plus_k_char_to_dl(35 downto 32);

LANE_STATE                 <= lane_state_from_lif;
RX_ERROR_CNT               <= rx_error_cnt_from_lif;
RX_ERROR_OVF               <= rx_error_ovf_from_lif;
LOSS_SIGNAL                <= no_signal_from_lcwd;
RX_POLARITY                <= invert_rx_bits_from_lif;
FAR_END_CAPA               <= far_end_capa_i;
lane_active_dl_i           <= enable_transm_data_from_lif;

QUAD0_rxp(0)               <= RX_POS;
QUAD0_rxn(0)               <= RX_NEG;
TX_POS                     <= QUAD0_txp(0);
TX_NEG                     <= QUAD0_txn(0);

RST_TX_DONE                <= INTF0_rst_tx_done_out_0;

end architecture rtl;
