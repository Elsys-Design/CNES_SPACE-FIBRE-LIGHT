// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_PHY_MS_DEFINES_VH
`else
`define B_HBM_PHY_MS_DEFINES_VH

// Look-up table parameters
//

`define HBM_PHY_MS_ADDR_N  43
`define HBM_PHY_MS_ADDR_SZ 32
`define HBM_PHY_MS_DATA_SZ 32

// Attribute addresses
//

`define HBM_PHY_MS__CFG0    32'h00000000
`define HBM_PHY_MS__CFG0_SZ 32

`define HBM_PHY_MS__CFG1    32'h00000001
`define HBM_PHY_MS__CFG1_SZ 29

`define HBM_PHY_MS__CFG10    32'h00000002
`define HBM_PHY_MS__CFG10_SZ 19

`define HBM_PHY_MS__CFG11    32'h00000003
`define HBM_PHY_MS__CFG11_SZ 11

`define HBM_PHY_MS__CFG12    32'h00000004
`define HBM_PHY_MS__CFG12_SZ 32

`define HBM_PHY_MS__CFG13    32'h00000005
`define HBM_PHY_MS__CFG13_SZ 16

`define HBM_PHY_MS__CFG14    32'h00000006
`define HBM_PHY_MS__CFG14_SZ 16

`define HBM_PHY_MS__CFG15    32'h00000007
`define HBM_PHY_MS__CFG15_SZ 28

`define HBM_PHY_MS__CFG16    32'h00000008
`define HBM_PHY_MS__CFG16_SZ 12

`define HBM_PHY_MS__CFG17    32'h00000009
`define HBM_PHY_MS__CFG17_SZ 16

`define HBM_PHY_MS__CFG18    32'h0000000a
`define HBM_PHY_MS__CFG18_SZ 32

`define HBM_PHY_MS__CFG19    32'h0000000b
`define HBM_PHY_MS__CFG19_SZ 32

`define HBM_PHY_MS__CFG2    32'h0000000c
`define HBM_PHY_MS__CFG2_SZ 32

`define HBM_PHY_MS__CFG20    32'h0000000d
`define HBM_PHY_MS__CFG20_SZ 32

`define HBM_PHY_MS__CFG21    32'h0000000e
`define HBM_PHY_MS__CFG21_SZ 16

`define HBM_PHY_MS__CFG22    32'h0000000f
`define HBM_PHY_MS__CFG22_SZ 3

`define HBM_PHY_MS__CFG23    32'h00000010
`define HBM_PHY_MS__CFG23_SZ 11

`define HBM_PHY_MS__CFG24    32'h00000011
`define HBM_PHY_MS__CFG24_SZ 14

`define HBM_PHY_MS__CFG25    32'h00000012
`define HBM_PHY_MS__CFG25_SZ 16

`define HBM_PHY_MS__CFG26    32'h00000013
`define HBM_PHY_MS__CFG26_SZ 12

`define HBM_PHY_MS__CFG27    32'h00000014
`define HBM_PHY_MS__CFG27_SZ 12

`define HBM_PHY_MS__CFG28    32'h00000015
`define HBM_PHY_MS__CFG28_SZ 12

`define HBM_PHY_MS__CFG29    32'h00000016
`define HBM_PHY_MS__CFG29_SZ 12

`define HBM_PHY_MS__CFG3    32'h00000017
`define HBM_PHY_MS__CFG3_SZ 21

`define HBM_PHY_MS__CFG31    32'h00000018
`define HBM_PHY_MS__CFG31_SZ 12

`define HBM_PHY_MS__CFG32    32'h00000019
`define HBM_PHY_MS__CFG32_SZ 16

`define HBM_PHY_MS__CFG33    32'h0000001a
`define HBM_PHY_MS__CFG33_SZ 4

`define HBM_PHY_MS__CFG34    32'h0000001b
`define HBM_PHY_MS__CFG34_SZ 16

`define HBM_PHY_MS__CFG35    32'h0000001c
`define HBM_PHY_MS__CFG35_SZ 16

`define HBM_PHY_MS__CFG36    32'h0000001d
`define HBM_PHY_MS__CFG36_SZ 16

`define HBM_PHY_MS__CFG37    32'h0000001e
`define HBM_PHY_MS__CFG37_SZ 16

`define HBM_PHY_MS__CFG38    32'h0000001f
`define HBM_PHY_MS__CFG38_SZ 9

`define HBM_PHY_MS__CFG39    32'h00000020
`define HBM_PHY_MS__CFG39_SZ 16

`define HBM_PHY_MS__CFG4    32'h00000021
`define HBM_PHY_MS__CFG4_SZ 9

`define HBM_PHY_MS__CFG40    32'h00000022
`define HBM_PHY_MS__CFG40_SZ 16

`define HBM_PHY_MS__CFG41    32'h00000023
`define HBM_PHY_MS__CFG41_SZ 18

`define HBM_PHY_MS__CFG42    32'h00000024
`define HBM_PHY_MS__CFG42_SZ 9

`define HBM_PHY_MS__CFG5    32'h00000025
`define HBM_PHY_MS__CFG5_SZ 8

`define HBM_PHY_MS__CFG6    32'h00000026
`define HBM_PHY_MS__CFG6_SZ 32

`define HBM_PHY_MS__CFG7    32'h00000027
`define HBM_PHY_MS__CFG7_SZ 16

`define HBM_PHY_MS__CFG8    32'h00000028
`define HBM_PHY_MS__CFG8_SZ 32

`define HBM_PHY_MS__CFG9    32'h00000029
`define HBM_PHY_MS__CFG9_SZ 32

`define HBM_PHY_MS__SIM_MODEL_TYPE    32'h0000002a
`define HBM_PHY_MS__SIM_MODEL_TYPE_SZ 24

`endif  // B_HBM_PHY_MS_DEFINES_VH