LIBRARY ieee ;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library work;
use work.pkg_simu.all;

entity tb_ppl_word_alignment is
end entity;

architecture tb of tb_ppl_word_alignment is

component ppl_64_word_alignment is
  port (
    RST_N                   : in  std_logic;                                          --! global reset
    CLK                     : in  std_logic;                                          --! Clock generated by HSSL IP
    -- ppm64_rx_sync_fsm (PLRSF) interface
    DATA_RX_PLWA            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! 64-bit data to lane_ctrl_word_detect
    VALID_K_CHARAC_PLWA     : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! 8-bit valid K character flags to lane_ctrl_word_detect
    DATA_RDY_PLWA           : out std_logic;                                          --! Data valid flag to lane_ctrl_word_detect
    INVALID_CHAR_PLWA       : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Invalid character flags from PLWA
    DISPARITY_ERR_PLWA      : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Disparity error flags from PLWA 
    RX_WORD_IS_ALIGNED_PLWA : out std_logic;                                          --! RX word is aligned from PLWA 
    COMMA_DET_PLWA          : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flag indicates that a comma is detected on the word receive from PLWA 
    -- HSSL IP interface
    DATA_RX_HSSL            : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! 64-bit data from HSSL IP
    VALID_K_CHARAC_HSSL     : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! 8-bit valid K character flags from HSSL IP
    INVALID_CHAR_HSSL       : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Invalid character flags from HSSL IP
    DISPARITY_ERR_HSSL      : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Disparity error flags from HSSL IP
    RX_WORD_IS_ALIGNED_HSSL : in  std_logic;                                          --! RX word is aligned from HSSL IP
    COMMA_DET_HSSL          : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0)  --! Flag indicates that a comma is detected on the word receive
   );
end component;



----------------------------- Stimulus signals
constant period                : time := 13.334 ns;
----- inputs
signal RST_N                   : std_logic                                          := '1';
signal CLK                     : std_logic                                          := '0';
signal DATA_RX_HSSL            : std_logic_vector(C_DATA_LENGTH-1 downto 0)         := (others =>'0');
signal VALID_K_CHARAC_HSSL     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0) := (others =>'0');
signal INVALID_CHAR_HSSL       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0):= (others => '0');
signal DISPARITY_ERR_HSSL      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0):= (others => '0');
signal RX_WORD_IS_ALIGNED_HSSL : std_logic                                          := '0';
signal COMMA_DET_HSSL          : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0) := (others=> '0');

----- Outputs
signal DATA_RX_PLWA            : std_logic_vector(C_DATA_LENGTH-1 downto 0);
signal VALID_K_CHARAC_PLWA     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
signal DATA_RDY_PLWA           : std_logic;
signal INVALID_CHAR_PLWA       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);
signal DISPARITY_ERR_PLWA      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);
signal RX_WORD_IS_ALIGNED_PLWA : std_logic;
signal COMMA_DET_PLWA          : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);

begin

-- Instantiate the DUT
DUT : ppl_64_word_alignment
  port map(
    RST_N                   => RST_N,
    CLK                     => CLK,
    DATA_RX_PLWA            => DATA_RX_PLWA,
    VALID_K_CHARAC_PLWA     => VALID_K_CHARAC_PLWA,
    DATA_RDY_PLWA           => DATA_RDY_PLWA,
    INVALID_CHAR_PLWA       => INVALID_CHAR_PLWA,
    DISPARITY_ERR_PLWA      => DISPARITY_ERR_PLWA,
    RX_WORD_IS_ALIGNED_PLWA => RX_WORD_IS_ALIGNED_PLWA,
    COMMA_DET_PLWA          => COMMA_DET_PLWA,
    DATA_RX_HSSL            => DATA_RX_HSSL,
    VALID_K_CHARAC_HSSL     => VALID_K_CHARAC_HSSL,
    INVALID_CHAR_HSSL       => INVALID_CHAR_HSSL, 
    DISPARITY_ERR_HSSL      => DISPARITY_ERR_HSSL,
    RX_WORD_IS_ALIGNED_HSSL => RX_WORD_IS_ALIGNED_HSSL,
    COMMA_DET_HSSL          => COMMA_DET_HSSL
  );

-- Clock generation process: 150 MHz clock
clk_gen : process
begin
  CLK <= not CLK;
  wait for period / 2;
end process;

-- Main stimulus process
scenario : process
  variable test_failed : boolean := false;
begin
  log_info("Applying reset");
  RST_N <= '0';
  wait for 10 us;
  wait until rising_edge(CLK);
  RST_N <= '1';
  wait for  1 us;
  -------------------------
  --     Start TEST      --
  -------------------------
  log_info("Star test");
  -------------------------
  -- Alignment on byte 0 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 0");
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  -- 2 words and a comma
  COMMA_DET_HSSL         <= "00000001";
  VALID_K_CHARAC_HSSL     <= "00000001";
  DATA_RX_HSSL           <= x"07060504030201BC";
  wait until rising_edge(CLK);
  -- new 2 words without comma
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0F0E0D0C0B0A0908";
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"0F0E0D0C0B0A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  wait until rising_edge(CLK);

  -------------------------
  -- Alignment on byte 1 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 1");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000010";
  VALID_K_CHARAC_HSSL     <= "00000010";
  DATA_RX_HSSL           <= x"060504030201BC99";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0E0D0C0B0A090807";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"000E0D0C0B0A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 2 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 2");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000100";
  VALID_K_CHARAC_HSSL     <= "00000100";
  DATA_RX_HSSL           <= x"0504030201BC9999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0D0C0B0A09080706";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"00000D0C0B0A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 3 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 3");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00001000";
  VALID_K_CHARAC_HSSL     <= "00001000";
  DATA_RX_HSSL           <= x"04030201BC999999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0C0B0A0908070605";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"0000000C0B0A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 4 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 4");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00010000";
  VALID_K_CHARAC_HSSL     <= "00010000";
  DATA_RX_HSSL           <= x"030201BC99999999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0B0A090807060504";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"000000000B0A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 5 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 5");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00100000";
  VALID_K_CHARAC_HSSL     <= "00100000";
  DATA_RX_HSSL           <= x"0201BC9999999999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0A09080706050403";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"00000000000A0908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 6 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 6");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "01000000";
  VALID_K_CHARAC_HSSL     <= "01000000";
  DATA_RX_HSSL           <= x"01BC999999999999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0908070605040302";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"0000000000000908", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  -------------------------
  -- Alignment on byte 7 --
  -------------------------
  report(LF & "##########################" & LF & "Alignment on byte 7");
  RX_WORD_IS_ALIGNED_HSSL <= '0';
  wait until rising_edge(CLK);
  RX_WORD_IS_ALIGNED_HSSL <= '1';
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "10000000";
  VALID_K_CHARAC_HSSL     <= "10000000";
  DATA_RX_HSSL           <= x"BC99999999999999";
  wait until rising_edge(CLK);
  COMMA_DET_HSSL         <= "00000000";
  VALID_K_CHARAC_HSSL     <= (others => '0');
  DATA_RX_HSSL           <= x"0807060504030201";
  wait until rising_edge(CLK);
  DATA_RX_HSSL           <= (others => '0');
  wait until rising_edge(CLK);
  -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"07060504030201BC", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000001"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
    -- check outputs
  check_equal("DATA_RX_PLWA"      ,  x"0000000000000008", DATA_RX_PLWA, test_failed);
  check_equal("VALID_K_CHARAC_PLWA", "00000000"         , VALID_K_CHARAC_PLWA, test_failed);
  wait until rising_edge(CLK);
  wait until rising_edge(CLK);

  -------------------------
  --       End TEST      --
  -------------------------

  log_info("All alignment tests completed.");
  wait for 1 us;
  log_test_result(test_failed);

  wait;
end process;

end tb;
