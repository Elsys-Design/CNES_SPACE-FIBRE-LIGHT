----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description :
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  
library phy_plus_lane_lib;
  use phy_plus_lane_lib.all;
  use phy_plus_lane_lib.pkg_phy_plus_lane.all;

entity lane_ctrl_word_insert is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP

      -- From DATA-LINK/TOP
      RD_DATA_FROM_DL                  : out std_logic;                       --! Read command to receive data from Data-link layer
      RD_DATA_VALID_FROM_DL            : in  std_logic;                       --! Data valid flag from Data-link layer
      CAPABILITY_FROM_DL               : in  std_logic_vector(07 downto 00);  --! Capability field from DATA-LINK layer
      DATA_TX_FROM_DL                  : in  std_logic_vector(31 downto 00);  --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_FROM_DL           : in  std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character from DATA-LINK layer
      NO_DATA_FROM_DL                  : in  std_logic;                       --! Flag to enable the send of IDLE words when no data should be available from Data-Link

      -- From/To skip_insertion
      WAIT_SEND_DATA_FROM_SKIP         : in  std_logic;                       --! Flag to indicates that the skip_insertion send a SKIP control word
      NEW_DATA_TO_SKIP                 : out std_logic;                       --! New data send to skip_insertion
      DATA_TX_TO_SKIP                  : out std_logic_vector(31 downto 00);  --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_TO_SKIP           : out std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character

      -- TX signals command from/to lane_init_fsm
      SEND_INIT1_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT2 control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD             : in  std_logic;                       --! Flag to send INIT3 control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA               : in  std_logic;                       --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS       : in  std_logic;                       --! Flag to send STANDBY control word x32
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  --! Standby reason from MIB
      SEND_32_LOSS_SIGNAL_CTRL_WORDS   : in  std_logic;                       --! Flag to send LOSS_SIGNAL control word x32
      LOST_CAUSE                       : in  std_logic_vector(01 downto 00);  --! Flag to indicate the reason of the LOST_SIGNAL
      STANDBY_SIGNAL_X32               : out std_logic;                       --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32                  : out std_logic                        --! Flag LOST_SIGNAL control word has been send x32
   );
end lane_ctrl_word_insert;

architecture rtl of lane_ctrl_word_insert is
----------------------------- Declaration signals -----------------------------

signal prbs_counter                 : unsigned(31 downto 00);                 --! PRBS value send during INIT1/2/3
signal init_word_sent               : std_logic;                              --! Indicates that the INIT1/2/3 control word has been send
signal send_stdby_cnt               : unsigned(04 downto 00);                 --! Standby counter x32
signal send_loss_sig_cnt            : unsigned(04 downto 00);                 --! Loss signal counter x32
signal no_data_from_dl_r            : std_logic;                              --! NO_DATA_FROM_DL with one clock cycle of delay
begin

-- Send data process
   p_send_data : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         RD_DATA_FROM_DL         <= '0';
         NEW_DATA_TO_SKIP        <= '0';
         DATA_TX_TO_SKIP         <= (others => '0');
         VALID_K_CHARAC_TO_SKIP  <= (others => '0');
         prbs_counter            <= (others => '0');
         init_word_sent          <= '0';
         send_stdby_cnt          <= (others => '0');
         STANDBY_SIGNAL_X32      <= '0';
         send_loss_sig_cnt       <= (others => '0');
         LOST_SIGNAL_X32         <= '0';
         no_data_from_dl_r       <= '0';

      elsif rising_edge(CLK) then

         no_data_from_dl_r <= NO_DATA_FROM_DL;

         if SEND_INIT1_CTRL_WORD = '1' or SEND_INIT2_CTRL_WORD = '1' or SEND_INIT3_CTRL_WORD = '1' then  -- When IP shall sent an INIT control word

            if prbs_counter = x"00000000" and init_word_sent = '0' then
               if SEND_INIT1_CTRL_WORD = '1' then                                                        -- When INIT1 control word shall be send
                  DATA_TX_TO_SKIP      <= C_INIT1_WORD;
               elsif SEND_INIT2_CTRL_WORD = '1' then                                                     -- When INIT2 control word shall be send
                  DATA_TX_TO_SKIP      <= C_INIT2_WORD;
               elsif SEND_INIT3_CTRL_WORD = '1' then                                                     -- When INIT3 control word shall be send
                  DATA_TX_TO_SKIP      <= CAPABILITY_FROM_DL & C_INIT3_WORD;
               end if;
               NEW_DATA_TO_SKIP        <= '1';
               VALID_K_CHARAC_TO_SKIP  <= x"1";                                                          -- Indicates that the Byte 1 is a K symbol
               init_word_sent          <= '1';                                                           -- Indicates that the first word have been sent
            elsif prbs_counter = C_PRBS_COUNTER_64 then
               prbs_counter            <= (others => '0');                                               -- Reset prbs counter
               NEW_DATA_TO_SKIP        <= '1';
               DATA_TX_TO_SKIP         <= std_logic_vector(prbs_counter);                                -- Send the 64th PRBS value
               VALID_K_CHARAC_TO_SKIP  <= x"0";                                                          -- Indicates no K symbol
               init_word_sent          <= '0';                                                           -- Reset flag
            elsif prbs_counter < C_PRBS_COUNTER_64 then
               prbs_counter            <= prbs_counter+1;                                                -- increment prbs counter by 1
               NEW_DATA_TO_SKIP        <= '1';
               DATA_TX_TO_SKIP         <= std_logic_vector(prbs_counter);                                -- Send 0 to 63 PRBS values
               VALID_K_CHARAC_TO_SKIP  <= x"0";                                                          -- Indicates no K symbol
            end if;


         elsif ENABLE_TRANSM_DATA = '1' then                                                             -- When the lane_init_fsm is in ACTIVE_ST
            NEW_DATA_TO_SKIP        <= '1';
            if ((no_data_from_dl_r = '0' and NO_DATA_FROM_DL = '1') or NO_DATA_FROM_DL = '0') and WAIT_SEND_DATA_FROM_SKIP = '0' then
               RD_DATA_FROM_DL         <= '1';
               if RD_DATA_VALID_FROM_DL ='1' then
                 DATA_TX_TO_SKIP         <= DATA_TX_FROM_DL;                                               -- Apply the data fornis by the DATA-LINK layer to the output
                 VALID_K_CHARAC_TO_SKIP  <= VALID_K_CHARAC_FROM_DL;                                        -- Indicates which byte is a K character from DATA-LINK layer
               else 
                  DATA_TX_TO_SKIP         <= C_IDLE_WORD;                                                   -- Sending IDLE control word
                  VALID_K_CHARAC_TO_SKIP  <= x"1";
               end if;
            elsif((no_data_from_dl_r = '0' and NO_DATA_FROM_DL = '1') or NO_DATA_FROM_DL = '0') and WAIT_SEND_DATA_FROM_SKIP = '1' then
               RD_DATA_FROM_DL         <= '0';
               if RD_DATA_VALID_FROM_DL ='1' then
                  DATA_TX_TO_SKIP         <= DATA_TX_FROM_DL;                                               -- Apply the data fornis by the DATA-LINK layer to the output
                  VALID_K_CHARAC_TO_SKIP  <= VALID_K_CHARAC_FROM_DL;                                        -- Indicates which byte is a K character from DATA-LINK layer
                else 
                   DATA_TX_TO_SKIP         <= C_IDLE_WORD;                                                   -- Sending IDLE control word
                   VALID_K_CHARAC_TO_SKIP  <= x"1";
                end if;
            else                                                         -- When no data has been send from DATA-LINK layer
               RD_DATA_FROM_DL         <= '1';
               DATA_TX_TO_SKIP         <= C_IDLE_WORD;                                                   -- Sending IDLE control word
               VALID_K_CHARAC_TO_SKIP  <= x"1";
            end if;


         elsif SEND_32_STANDBY_CTRL_WORDS = '1' then                                                     -- When the lane_init_fsm is in PREPARE_STANDBY_ST

            if send_stdby_cnt >= C_X32_SIGNAL then                                                       -- When 32 STANDBY control words has been send
               STANDBY_SIGNAL_X32      <= '1';                                                           -- Indicates to lane_init_fsm that the STANDBY control word x32 has been send                                                 -- Reset counter
            elsif send_stdby_cnt < C_X32_SIGNAL then                                                     -- else
               STANDBY_SIGNAL_X32      <= '0';                                                           -- Indicates to lane_init_fsm that the STANDBY control word x32 has not been send
               send_stdby_cnt          <= send_stdby_cnt+1;                                              -- Increment counter by 1
               NEW_DATA_TO_SKIP        <= '1';
               DATA_TX_TO_SKIP         <= STANDBY_REASON & C_STANDBY_WORD;                               -- Send STANDBY control word
               VALID_K_CHARAC_TO_SKIP  <= x"1";                                                          -- Indicates that the Byte 1 is a K symbol
            end if;


         elsif SEND_32_LOSS_SIGNAL_CTRL_WORDS = '1' then                                                 -- When the lane_init_fsm is in LOSS_OF_SIGNAL_ST

            if send_loss_sig_cnt >= C_X32_SIGNAL then                                                    -- When 32 LOSS_SIGNAL control words has been send
               LOST_SIGNAL_X32         <= '1';                                                           -- Indicates to lane_init_fsm that the LOSS_SIGNAL control word x32 has been send
            elsif send_loss_sig_cnt < C_X32_SIGNAL then                                                  -- else
               LOST_SIGNAL_X32         <= '0';                                                           -- Indicates to lane_init_fsm that the LOSS_SIGNAL control word x32 has not been send
               send_loss_sig_cnt       <= send_loss_sig_cnt+1;                                           -- Increment counter by 1
               NEW_DATA_TO_SKIP        <= '1';
               DATA_TX_TO_SKIP         <= "000000" & LOST_CAUSE & C_LOST_SIG_WORD;                        -- Send LOSS_SIGNAL control word
               VALID_K_CHARAC_TO_SKIP  <= x"1";                                                          -- Indicates that the Byte 1 is a K symbol
            end if;

         else
            RD_DATA_FROM_DL         <= '0';
            NEW_DATA_TO_SKIP        <= '0';
            DATA_TX_TO_SKIP         <= (others => '0');                                                  -- Reset all counters and flags
            VALID_K_CHARAC_TO_SKIP  <= (others => '0');
            prbs_counter            <= (others => '0');
            init_word_sent          <= '0';
            send_stdby_cnt          <= (others => '0');
            STANDBY_SIGNAL_X32      <= '0';
            send_loss_sig_cnt       <= (others => '0');
            LOST_SIGNAL_X32         <= '0';
         end if;

      end if;
   end process p_send_data;

end architecture rtl;
