-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibre_Light Versal target
--
-- Creation date : 03/09/2024
--
-- Description : This module implement the Physical and Lane layer of an IP
-- SpaceFibre Light.
-- The Physical layer is carried by an Xilinx IP
-- The Lane layer is carried by owner's code and an Xilinx IP
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library unisim;
use unisim.vcomponents.all;

library commun;
use commun.all;

entity phy_plus_lane_64b_to_32b is
   port(
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Main clock
      -- Reset_gen interface 
      LANE_RESET_PPL_OUT               : out std_logic;
      RST_TXCLK_N                      : in  std_logic;                       --! Synchronous reset on clock generated by GTY PLL
      CLK_TX_OUT                       : out std_logic;                       --! Clock generated by manufacturer IP
      RST_TX_DONE                      : out std_logic;                       --! Up when internal rx reset done
      -- CLK GTY signals
      CLK_GTY                          : in std_logic;                        --! Clock for the extended phy layer IP
      -- FROM Data-link layer
      DATA_TX                          : in  std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be send from Data-Link Layer
      LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer
      CAPABILITY_TX                    : in  std_logic_vector(07 downto 00);  --! Capability field send in INIT3 control word
      NEW_DATA_TX                      : in  std_logic;                       --! Flag new data
      VALID_K_CHARAC_TX                : in  std_logic_vector(03 downto 00);  --! 4-bit valid K character flags from Data-link layer
      FIFO_TX_FULL                     : out std_logic;                       --! FiFo TX full flag

      -- TO Data-link layer
      FIFO_RX_RD_EN                    : in  std_logic;                       --! FiFo RX read enable flag
      DATA_RX                          : out std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be received to Data-Link Layer
      FIFO_RX_EMPTY                    : out std_logic;                       --! FiFo RX empty flag
      FIFO_RX_DATA_VALID               : out std_logic;                       --! FiFo RX data valid flag
      VALID_K_CHARAC_RX                : out std_logic_vector(03 downto 00);  --! 4-bit valid K character flags to Data-link layer
      FAR_END_CAPA_DL                  : out std_logic_vector(07 downto 00);  --! Capability field receive in INIT3 control word
      LANE_ACTIVE_DL                   : out std_logic;                       --! Lane Active flag for the DATA Link Layer

      -- FROM/TO Outside
      TX_POS                           : out std_logic;                       --! Positive LVDS serial data send
      TX_NEG                           : out std_logic;                       --! Negative LVDS serial data send
      RX_POS                           : in  std_logic;                       --! Positive LVDS serial data received
      RX_NEG                           : in  std_logic;                       --! Negative LVDS serial data received

      -- PARAMETERS and STATUS
      LANE_START                       : in  std_logic;                       --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                       --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                       --! Asserts or de-asserts LaneReset for the lane
      PARALLEL_LOOPBACK_EN             : in  std_logic;                       --! Enables or disables the parallel loopback for the lane
      STANDBY_REASON_MIB                   : in  std_logic_vector(07 downto 00);  --! In case of error, pauses communication
      NEAR_END_SERIAL_LB_EN            : in  std_logic;                       --! Enables or disables the near-end serial loopback for the lane
      FAR_END_SERIAL_LB_EN             : in  std_logic;                       --! Enables or disables the far-end serial loopback for the lane

      LANE_STATE                       : out std_logic_vector(03 downto 00);  --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic;                       --! Overflow flag of the RX_ERROR_CNT
      LOSS_SIGNAL                      : out std_logic;                       --! Set when no signal is received on RX link
      FAR_END_CAPA                     : out std_logic_vector(07 downto 00);  --! Capabilities field (INT3 flags)
      RX_POLARITY                      : out std_logic                        --! Set when the receiver polarity is inverted
   );
end phy_plus_lane_64b_to_32b;

architecture rtl of phy_plus_lane_64b_to_32b is
   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Modules Declaration -----------------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
   

   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Internal signals declaration --------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------

begin
   ------------------------------------------------------------------------------
   -- Instance of rx_sync_fsm module
   ------------------------------------------------------------------------------
   inst_rx_sync_fsm : rx_sync_fsm
   port map(
      CLK_SYS                          => CLK,
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- FROM Data-link layer
      LANE_RESET_DL                    => lane_reset_dl_i,
      -- TO lane_ctrl_word_detection
      DATA_RX_PLRSF                 => data_rx_from_rsf,
      VALID_K_CHARAC_PLRSF           => valid_k_charac_from_rsf,
      DATA_RDY_PLRSF                => data_rdy_from_rsf,
      -- FROM MANUFACTURER IP
      DATA_RX_HSSL                  => INTF0_RX0_ch_rxdata(31 downto 00),
      VALID_K_CHARAC_HSSL            => INTF0_RX0_ch_rxctrl0(03 downto 00),
      DATA_RDY_HSSL                 => INTF0_RX0_ch_rxdatavalid(0),
      INVALID_CHAR_HSSL             => INTF0_RX0_ch_rxctrl3(03 downto 00),
      DISPARITY_ERR_HSSL            => INTF0_RX0_ch_rxctrl1(03 downto 00),
      RX_WORD_REALIGN_HSSL          => INTF0_RX0_ch_rxbyterealign(0),
      COMMA_DET_HSSL                => INTF0_RX0_ch_rxctrl2(0),
      -- PARAMETERS
      LANE_RESET                       => LANE_RESET
   );
   ------------------------------------------------------------------------------
   -- Instance of TX BufG_GT_wrapper module for TX clock
   ------------------------------------------------------------------------------
      inst_bufg_gt_tx_clock : BufG_GT_bd_wrapper
         port map(
           gt_bufgtce_0                   => '1',
           gt_bufgtcemask_0               => '0',
           gt_bufgtclr_0                  => '0',
           gt_bufgtclrmask_0              => '0',
           gt_bufgtdiv_0                  => "000",
           outclk_0                       => QUAD0_TX0_outclk,
           usrclk_0                       => clk_tx
         );

   reset <= not RST_N or LANE_RESET or lane_reset_dl_i;

   -- Near-End and Far-End loopback drivin function
   QUAD0_ch0_loopback         <= "010"    when NEAR_END_SERIAL_LB_EN = '1' else
                                 "100"    when FAR_END_SERIAL_LB_EN = '1'  else
                                 "000";

   -- Clock Data recovery drivin function
   INTF0_RX0_ch_rxcdrhold     <= "0"      when cdr_from_lif = '1' else "1";
   INTF0_RX0_ch_rxcdrovrden   <= "0"      when cdr_from_lif = '1' else "0";

   -- Disable transmitter and/or receiver drinvin function
   INTF0_TX0_ch_txpd          <= "11"     when transmitter_dis_from_lif = '1' else "00";
   INTF0_RX0_ch_rxpd          <= "11"     when receiver_dis_from_lif = '1' else "00";

   ------------------------------------------------------------------------------
   -- Instance of extended_phy_layer module
   ------------------------------------------------------------------------------
  inst_extended_phy_layer_wrapper : extended_phy_layer_wrapper
   port map(
     INTF0_RX0_ch_rxbufstatus_0           => open,
     INTF0_RX0_ch_rxbyteisaligned_0       => open,
     INTF0_RX0_ch_rxbyterealign_0         => INTF0_RX0_ch_rxbyterealign,
     INTF0_RX0_ch_rxcdrhold_0             => INTF0_RX0_ch_rxcdrhold,
     INTF0_RX0_ch_rxcdrovrden_0           => INTF0_RX0_ch_rxcdrovrden,
     INTF0_RX0_ch_rxcomsasdet_0           => open,
     INTF0_RX0_ch_rxctrl0_0               => INTF0_RX0_ch_rxctrl0,
     INTF0_RX0_ch_rxctrl1_0               => INTF0_RX0_ch_rxctrl1,
     INTF0_RX0_ch_rxctrl2_0               => INTF0_RX0_ch_rxctrl2,
     INTF0_RX0_ch_rxctrl3_0               => INTF0_RX0_ch_rxctrl3,
     INTF0_RX0_ch_rxdata_0                => INTF0_RX0_ch_rxdata,
     INTF0_RX0_ch_rxdatavalid_0           => INTF0_RX0_ch_rxdatavalid,
     INTF0_RX0_ch_rxpd_0                  => INTF0_RX0_ch_rxpd,
     INTF0_RX0_ch_rxpolarity_0(0)         => invert_rx_bits_from_lif,
     INTF0_RX0_ch_rxrate_0                => "00000000",
     INTF0_RX_clr_out_0                   => open,
     INTF0_RX_clrb_leaf_out_0             => open,
     INTF0_TX0_ch_txbufstatus_0           => open,
     INTF0_TX0_ch_txctrl0_0               => "0000000000000000",
     INTF0_TX0_ch_txctrl1_0               => "0000000000000000",
     INTF0_TX0_ch_txctrl2_0               => valid_k_charac_from_si,
     INTF0_TX0_ch_txdata                  => data_tx_from_si,
     INTF0_TX0_ch_txpd_0                  => INTF0_TX0_ch_txpd,
     INTF0_TX0_ch_txrate_0                => "00000000",
     INTF0_TX_clr_out_0                   => open,
     INTF0_TX_clrb_leaf_out_0             => open,
     INTF0_rst_all_in_0                   => reset,
     INTF0_rst_rx_datapath_in_0           => '0',
     INTF0_rst_rx_done_out_0              => open,
     INTF0_rst_rx_pll_and_datapath_in_0   => '0',
     INTF0_rst_tx_datapath_in_0           => '0',
     INTF0_rst_tx_done_out_0              => INTF0_rst_tx_done_out_0,
     INTF0_rst_tx_pll_and_datapath_in_0   => '0',
     QUAD0_GTREFCLK0_0                    => CLK_GTY,
     QUAD0_GT_DEBUG_0_gpi                 => x"00000000",
     QUAD0_GT_DEBUG_0_gpo                 => open,
     QUAD0_RX0_outclk_0                   => open,
     QUAD0_RX0_usrclk_0                   => clk_tx,--QUAD0_TX0_outclk,
     QUAD0_TX0_outclk_0                   => QUAD0_TX0_outclk,
     QUAD0_TX0_usrclk_0                   => clk_tx, --QUAD0_TX0_outclk,
     QUAD0_hsclk0_lcplllock_0             => QUAD0_hsclk0_lcplllock,
     Quad0_CH0_DEBUG_0_ch_loopback        => QUAD0_ch0_loopback,
     Quad0_GT_Serial_0_grx_n              => QUAD0_rxn,
     Quad0_GT_Serial_0_grx_p              => QUAD0_rxp,
     Quad0_GT_Serial_0_gtx_n              => QUAD0_txn,
     Quad0_GT_Serial_0_gtx_p              => QUAD0_txp,
     gtpowergood_0                        => open,
     gtwiz_freerun_clk_0                  => CLK
   );

inst_spacefibre_hssl_64b: SpaceFibre_64b
port map (
    -- Serial ports
    hssl_clock_i            => hssl_tx_clock_i,
    rx0n                    => lane_rx_rx0n,
    rx0p                    => lane_rx_rx0p,
    rx1n                    => '1',
    rx1p                    => '0',
    rx2n                    => '1',
    rx2p                    => '0',
    rx3n                    => '1',
    rx3p                    => '0',
    tx0n                    => lane_tx_tx0n,
    tx0p                    => lane_tx_tx0p,
    tx1n                    => open,
    tx1p                    => open,
    tx2n                    => open,
    tx2p                    => open,
    tx3n                    => open,
    tx3p                    => open,
    -- Clocks
    ckrefn                  => ckrefn,
    ckrefp                  => ckrefp,
    clock_o                 => CLK_HSSL,
    -- PMA PLL ports (do not touch)
    dyn_cfg_en_i            => '1',
    dyn_addr_i              => "0000",
    dyn_calibration_cs_n_i  => '1',
    dyn_lane_cs_n_i         => "1111",
    dyn_wdata_i             => "000000000000",
    dyn_wdata_sel_i         => '0',
    dyn_we_n_i              => '1',
    -- PMA PLL ports
    pll_pma_lock_analog     => pll_pma_lock_analog_tx,
    pll_pma_pwr_up_i        => pll_pma_pwr_up_tx,
    pll_pma_rst_n_i         => pll_pma_rst_n_tx,
    pll_lock                => open,
    -- TX ports
    tx0_busy_o              => tx_busy,
    tx0_clk_ena_i           => TX_CLK_ENA,
    tx0_clk_o               => TX_CLK_HSSL,
    tx0_data_i              => tx_data,
    tx0_ctrl_driver_pwrdwn_n_i => tx_driver_pwrdwn_n,
    tx0_rst_n_i             => tx_rst_n,
    tx0_ctrl_char_is_k_i    => tx_ctrl_char_is_k,
    -- RX ports
    rx0_busy_o              => open,
    rx0_ctrl_el_buff_stat_o => open,
    rx0_ctrl_char_is_aligned_o => open,
    rx0_ctrl_char_is_comma_o => open,
    rx0_ctrl_char_is_f_o    => open,
    rx0_ctrl_char_is_k_o    => open,
    rx0_ctrl_disp_err_o     => open,
    rx0_ctrl_not_in_table_o => open,
    rx0_ctrl_valid_realign_o => open,
    rx0_data_o              => open,
    rx0_ovs_bit_sel_i       => "00",
    rx0_eye_rst_i           => '0',
    rx0_pma_ll_fast_locked_o => open,
    rx0_pma_ll_slow_locked_o => rx_pma_ll_slow_locked,
    rx0_pma_loss_of_signal_o => RX_PMA_LOSS_OF_SIGNAL_HSSL,
    rx0_pma_pll_lock_o      => open,
    rx0_pma_pll_lock_track_o => open,
    rx0_pma_rst_n_i         => rx_pma_rst_n,
    rx0_pma_pwr_up_i        => rx_pma_pwr_up,
    rx0_rst_n_i             => rx_rst_n,
    rx0_test_o              => open,
    rx0_replace_en_i        => '0',
    rx0_align_sync_i        => rx_align_sync,
    rx0_el_buff_rst_i       => '0'
);


  -- Inputs/Outputs
CLK_TX_OUT                 <= clk_tx;

data_plus_k_char_from_dl   <= VALID_K_CHARAC_TX & DATA_TX;
DATA_RX                    <= data_plus_k_char_to_dl(31 downto 00);
VALID_K_CHARAC_RX          <= data_plus_k_char_to_dl(35 downto 32);

LANE_STATE                 <= lane_state_from_lif;
RX_ERROR_CNT               <= rx_error_cnt_from_lif;
RX_ERROR_OVF               <= rx_error_ovf_from_lif;
LOSS_SIGNAL                <= no_signal_from_lcwd;
RX_POLARITY                <= invert_rx_bits_from_lif;
FAR_END_CAPA               <= far_end_capa_i;
lane_active_dl_i           <= ENABLE_TRANSM_DATA_PLIF_from_lif;

QUAD0_rxp(0)               <= RX_POS;
QUAD0_rxn(0)               <= RX_NEG;
TX_POS                     <= QUAD0_txp(0);
TX_NEG                     <= QUAD0_txn(0);

RST_TX_DONE                <= INTF0_rst_tx_done_out_0;

end architecture rtl;
