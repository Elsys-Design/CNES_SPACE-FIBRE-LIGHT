`include "B_DFE_PRACH_defines.vh"

reg [`DFE_PRACH_DATA_SZ-1:0] ATTR [0:`DFE_PRACH_ADDR_N-1];
real ACTIVE_DUTYCYCLE_REG = ACTIVE_DUTYCYCLE;
real CLK_FREQ_REG = CLK_FREQ;
real DECIMATION_RATE_REG = DECIMATION_RATE;
real INCOMING_SAMPLE_RATE_REG = INCOMING_SAMPLE_RATE;
reg [`DFE_PRACH__INCOMING_SAMPLE_RATE_STR_SZ:1] INCOMING_SAMPLE_RATE_STR_REG = INCOMING_SAMPLE_RATE_STR;
real NUM_ACTIVE_ANTENNAS_REG = NUM_ACTIVE_ANTENNAS;
real NUM_ACTIVE_CHANNELS_REG = NUM_ACTIVE_CHANNELS;
reg [`DFE_PRACH__XPA_CFG0_SZ-1:0] XPA_CFG0_REG = XPA_CFG0;

initial begin
  ATTR[`DFE_PRACH__ACTIVE_DUTYCYCLE] = $realtobits(ACTIVE_DUTYCYCLE);
  ATTR[`DFE_PRACH__CLK_FREQ] = $realtobits(CLK_FREQ);
  ATTR[`DFE_PRACH__DECIMATION_RATE] = $realtobits(DECIMATION_RATE);
  ATTR[`DFE_PRACH__INCOMING_SAMPLE_RATE] = $realtobits(INCOMING_SAMPLE_RATE);
  ATTR[`DFE_PRACH__INCOMING_SAMPLE_RATE_STR] = INCOMING_SAMPLE_RATE_STR;
  ATTR[`DFE_PRACH__NUM_ACTIVE_ANTENNAS] = $realtobits(NUM_ACTIVE_ANTENNAS);
  ATTR[`DFE_PRACH__NUM_ACTIVE_CHANNELS] = $realtobits(NUM_ACTIVE_CHANNELS);
  ATTR[`DFE_PRACH__XPA_CFG0] = XPA_CFG0;
end

always @(trig_attr) begin
  ACTIVE_DUTYCYCLE_REG = $bitstoreal(ATTR[`DFE_PRACH__ACTIVE_DUTYCYCLE]);
  CLK_FREQ_REG = $bitstoreal(ATTR[`DFE_PRACH__CLK_FREQ]);
  DECIMATION_RATE_REG = $bitstoreal(ATTR[`DFE_PRACH__DECIMATION_RATE]);
  INCOMING_SAMPLE_RATE_REG = $bitstoreal(ATTR[`DFE_PRACH__INCOMING_SAMPLE_RATE]);
  INCOMING_SAMPLE_RATE_STR_REG = ATTR[`DFE_PRACH__INCOMING_SAMPLE_RATE_STR];
  NUM_ACTIVE_ANTENNAS_REG = $bitstoreal(ATTR[`DFE_PRACH__NUM_ACTIVE_ANTENNAS]);
  NUM_ACTIVE_CHANNELS_REG = $bitstoreal(ATTR[`DFE_PRACH__NUM_ACTIVE_CHANNELS]);
  XPA_CFG0_REG = ATTR[`DFE_PRACH__XPA_CFG0];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DFE_PRACH_ADDR_SZ-1:0] addr;
  input  [`DFE_PRACH_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DFE_PRACH_DATA_SZ-1:0] read_attr;
  input  [`DFE_PRACH_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
