`include "B_DSP_FP_INREG_defines.vh"

reg [`DSP_FP_INREG_DATA_SZ-1:0] ATTR [0:`DSP_FP_INREG_ADDR_N-1];
reg [`DSP_FP_INREG__ACASCREG_SZ-1:0] ACASCREG_REG = ACASCREG;
reg [`DSP_FP_INREG__AREG_SZ-1:0] AREG_REG = AREG;
reg [`DSP_FP_INREG__A_FPTYPE_SZ:1] A_FPTYPE_REG = A_FPTYPE;
reg [`DSP_FP_INREG__A_INPUT_SZ:1] A_INPUT_REG = A_INPUT;
reg [`DSP_FP_INREG__BCASCSEL_SZ:1] BCASCSEL_REG = BCASCSEL;
reg [`DSP_FP_INREG__B_D_FPTYPE_SZ:1] B_D_FPTYPE_REG = B_D_FPTYPE;
reg [`DSP_FP_INREG__B_INPUT_SZ:1] B_INPUT_REG = B_INPUT;
reg [`DSP_FP_INREG__FPBREG_SZ-1:0] FPBREG_REG = FPBREG;
reg [`DSP_FP_INREG__FPDREG_SZ-1:0] FPDREG_REG = FPDREG;
reg IS_RSTA_INVERTED_REG = IS_RSTA_INVERTED;
reg IS_RSTB_INVERTED_REG = IS_RSTB_INVERTED;
reg [`DSP_FP_INREG__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;

initial begin
  ATTR[`DSP_FP_INREG__ACASCREG] = ACASCREG;
  ATTR[`DSP_FP_INREG__AREG] = AREG;
  ATTR[`DSP_FP_INREG__A_FPTYPE] = A_FPTYPE;
  ATTR[`DSP_FP_INREG__A_INPUT] = A_INPUT;
  ATTR[`DSP_FP_INREG__BCASCSEL] = BCASCSEL;
  ATTR[`DSP_FP_INREG__B_D_FPTYPE] = B_D_FPTYPE;
  ATTR[`DSP_FP_INREG__B_INPUT] = B_INPUT;
  ATTR[`DSP_FP_INREG__FPBREG] = FPBREG;
  ATTR[`DSP_FP_INREG__FPDREG] = FPDREG;
  ATTR[`DSP_FP_INREG__IS_RSTA_INVERTED] = IS_RSTA_INVERTED;
  ATTR[`DSP_FP_INREG__IS_RSTB_INVERTED] = IS_RSTB_INVERTED;
  ATTR[`DSP_FP_INREG__RESET_MODE] = RESET_MODE;
end

always @(trig_attr) begin
  ACASCREG_REG = ATTR[`DSP_FP_INREG__ACASCREG];
  AREG_REG = ATTR[`DSP_FP_INREG__AREG];
  A_FPTYPE_REG = ATTR[`DSP_FP_INREG__A_FPTYPE];
  A_INPUT_REG = ATTR[`DSP_FP_INREG__A_INPUT];
  BCASCSEL_REG = ATTR[`DSP_FP_INREG__BCASCSEL];
  B_D_FPTYPE_REG = ATTR[`DSP_FP_INREG__B_D_FPTYPE];
  B_INPUT_REG = ATTR[`DSP_FP_INREG__B_INPUT];
  FPBREG_REG = ATTR[`DSP_FP_INREG__FPBREG];
  FPDREG_REG = ATTR[`DSP_FP_INREG__FPDREG];
  IS_RSTA_INVERTED_REG = ATTR[`DSP_FP_INREG__IS_RSTA_INVERTED];
  IS_RSTB_INVERTED_REG = ATTR[`DSP_FP_INREG__IS_RSTB_INVERTED];
  RESET_MODE_REG = ATTR[`DSP_FP_INREG__RESET_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FP_INREG_ADDR_SZ-1:0] addr;
  input  [`DSP_FP_INREG_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FP_INREG_DATA_SZ-1:0] read_attr;
  input  [`DSP_FP_INREG_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
