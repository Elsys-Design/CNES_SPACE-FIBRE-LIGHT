`include "B_DSP_FPA_OPM_REG_defines.vh"

reg [`DSP_FPA_OPM_REG_DATA_SZ-1:0] ATTR [0:`DSP_FPA_OPM_REG_ADDR_N-1];
reg [`DSP_FPA_OPM_REG__FPMPIPEREG_SZ-1:0] FPMPIPEREG_REG = FPMPIPEREG;
reg [`DSP_FPA_OPM_REG__FPOPMREG_SZ-1:0] FPOPMREG_REG = FPOPMREG;
reg [`DSP_FPA_OPM_REG__IS_FPOPMODE_INVERTED_SZ-1:0] IS_FPOPMODE_INVERTED_REG = IS_FPOPMODE_INVERTED;
reg IS_RSTFPOPMODE_INVERTED_REG = IS_RSTFPOPMODE_INVERTED;
reg [`DSP_FPA_OPM_REG__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;
reg [`DSP_FPA_OPM_REG__USE_MULT_SZ:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_FPA_OPM_REG__FPMPIPEREG] = FPMPIPEREG;
  ATTR[`DSP_FPA_OPM_REG__FPOPMREG] = FPOPMREG;
  ATTR[`DSP_FPA_OPM_REG__IS_FPOPMODE_INVERTED] = IS_FPOPMODE_INVERTED;
  ATTR[`DSP_FPA_OPM_REG__IS_RSTFPOPMODE_INVERTED] = IS_RSTFPOPMODE_INVERTED;
  ATTR[`DSP_FPA_OPM_REG__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_FPA_OPM_REG__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  FPMPIPEREG_REG = ATTR[`DSP_FPA_OPM_REG__FPMPIPEREG];
  FPOPMREG_REG = ATTR[`DSP_FPA_OPM_REG__FPOPMREG];
  IS_FPOPMODE_INVERTED_REG = ATTR[`DSP_FPA_OPM_REG__IS_FPOPMODE_INVERTED];
  IS_RSTFPOPMODE_INVERTED_REG = ATTR[`DSP_FPA_OPM_REG__IS_RSTFPOPMODE_INVERTED];
  RESET_MODE_REG = ATTR[`DSP_FPA_OPM_REG__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_FPA_OPM_REG__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FPA_OPM_REG_ADDR_SZ-1:0] addr;
  input  [`DSP_FPA_OPM_REG_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FPA_OPM_REG_DATA_SZ-1:0] read_attr;
  input  [`DSP_FPA_OPM_REG_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
