// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC_NIDB_DEFINES_VH
`else
`define B_NOC_NIDB_DEFINES_VH

// Look-up table parameters
//

`define NOC_NIDB_ADDR_N  30
`define NOC_NIDB_ADDR_SZ 32
`define NOC_NIDB_DATA_SZ 32

// Attribute addresses
//

`define NOC_NIDB__REG_ADDR_REMAP0    32'h00000000
`define NOC_NIDB__REG_ADDR_REMAP0_SZ 32

`define NOC_NIDB__REG_ADDR_REMAP1    32'h00000001
`define NOC_NIDB__REG_ADDR_REMAP1_SZ 16

`define NOC_NIDB__REG_ADDR_REMAP_MASK0    32'h00000002
`define NOC_NIDB__REG_ADDR_REMAP_MASK0_SZ 32

`define NOC_NIDB__REG_ADDR_REMAP_MASK1    32'h00000003
`define NOC_NIDB__REG_ADDR_REMAP_MASK1_SZ 16

`define NOC_NIDB__REG_BYPASS_CNTL    32'h00000004
`define NOC_NIDB__REG_BYPASS_CNTL_SZ 2

`define NOC_NIDB__REG_DCC_CNTR    32'h00000005
`define NOC_NIDB__REG_DCC_CNTR_SZ 10

`define NOC_NIDB__REG_ECC_CHK_EN    32'h00000006
`define NOC_NIDB__REG_ECC_CHK_EN_SZ 2

`define NOC_NIDB__REG_ERR_PKT_DROP_DIS    32'h00000007
`define NOC_NIDB__REG_ERR_PKT_DROP_DIS_SZ 3

`define NOC_NIDB__REG_IO_CHAR_EN    32'h00000008
`define NOC_NIDB__REG_IO_CHAR_EN_SZ 11

`define NOC_NIDB__REG_IO_CHAR_OUTPUT_MUX_SEL    32'h00000009
`define NOC_NIDB__REG_IO_CHAR_OUTPUT_MUX_SEL_SZ 11

`define NOC_NIDB__REG_IO_CNTRL    32'h0000000a
`define NOC_NIDB__REG_IO_CNTRL_SZ 11

`define NOC_NIDB__REG_LOOPBACK_CNTL    32'h0000000b
`define NOC_NIDB__REG_LOOPBACK_CNTL_SZ 3

`define NOC_NIDB__REG_NOC_CTL    32'h0000000c
`define NOC_NIDB__REG_NOC_CTL_SZ 16

`define NOC_NIDB__REG_P0_0_VCA_TOKEN    32'h0000000d
`define NOC_NIDB__REG_P0_0_VCA_TOKEN_SZ 32

`define NOC_NIDB__REG_P0_1_VCA_TOKEN    32'h0000000e
`define NOC_NIDB__REG_P0_1_VCA_TOKEN_SZ 32

`define NOC_NIDB__REG_RX_DELAY_EN    32'h0000000f
`define NOC_NIDB__REG_RX_DELAY_EN_SZ 10

`define NOC_NIDB__REG_RX_DW0_DELAY    32'h00000010
`define NOC_NIDB__REG_RX_DW0_DELAY_SZ 18

`define NOC_NIDB__REG_RX_DW1_DELAY    32'h00000011
`define NOC_NIDB__REG_RX_DW1_DELAY_SZ 18

`define NOC_NIDB__REG_RX_DW2_DELAY    32'h00000012
`define NOC_NIDB__REG_RX_DW2_DELAY_SZ 18

`define NOC_NIDB__REG_RX_DW3_DELAY    32'h00000013
`define NOC_NIDB__REG_RX_DW3_DELAY_SZ 18

`define NOC_NIDB__REG_RX_DW4_DELAY    32'h00000014
`define NOC_NIDB__REG_RX_DW4_DELAY_SZ 18

`define NOC_NIDB__REG_TX_DCC_DELAY    32'h00000015
`define NOC_NIDB__REG_TX_DCC_DELAY_SZ 8

`define NOC_NIDB__REG_VC0_ARPROT_SEL    32'h00000016
`define NOC_NIDB__REG_VC0_ARPROT_SEL_SZ 6

`define NOC_NIDB__REG_VC0_SMID_SEL    32'h00000017
`define NOC_NIDB__REG_VC0_SMID_SEL_SZ 20

`define NOC_NIDB__REG_VC1_AWPROT_SEL    32'h00000018
`define NOC_NIDB__REG_VC1_AWPROT_SEL_SZ 6

`define NOC_NIDB__REG_VC1_SMID_SEL    32'h00000019
`define NOC_NIDB__REG_VC1_SMID_SEL_SZ 20

`define NOC_NIDB__REG_VC4_ARPROT_SEL    32'h0000001a
`define NOC_NIDB__REG_VC4_ARPROT_SEL_SZ 6

`define NOC_NIDB__REG_VC4_SMID_SEL    32'h0000001b
`define NOC_NIDB__REG_VC4_SMID_SEL_SZ 20

`define NOC_NIDB__REG_VC5_AWPROT_SEL    32'h0000001c
`define NOC_NIDB__REG_VC5_AWPROT_SEL_SZ 6

`define NOC_NIDB__REG_VC5_SMID_SEL    32'h0000001d
`define NOC_NIDB__REG_VC5_SMID_SEL_SZ 20

`endif  // B_NOC_NIDB_DEFINES_VH