// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DCMAC_DEFINES_VH
`else
`define B_DCMAC_DEFINES_VH

// Look-up table parameters
//

`define DCMAC_ADDR_N  1254
`define DCMAC_ADDR_SZ 32
`define DCMAC_DATA_SZ 64

// Attribute addresses
//

`define DCMAC__C0_CTL_PCS_RX_TS_EN    32'h00000000
`define DCMAC__C0_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_ACK    32'h00000001
`define DCMAC__C0_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_ETYPE_GCP    32'h00000002
`define DCMAC__C0_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_ETYPE_GPP    32'h00000003
`define DCMAC__C0_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_ETYPE_PCP    32'h00000004
`define DCMAC__C0_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_ETYPE_PPP    32'h00000005
`define DCMAC__C0_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_MCAST_GCP    32'h00000006
`define DCMAC__C0_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_MCAST_GPP    32'h00000007
`define DCMAC__C0_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_MCAST_PCP    32'h00000008
`define DCMAC__C0_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_MCAST_PPP    32'h00000009
`define DCMAC__C0_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_OPCODE_GCP    32'h0000000a
`define DCMAC__C0_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_OPCODE_GPP    32'h0000000b
`define DCMAC__C0_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_OPCODE_PCP    32'h0000000c
`define DCMAC__C0_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_OPCODE_PPP    32'h0000000d
`define DCMAC__C0_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_PREAMBLE    32'h0000000e
`define DCMAC__C0_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_SA_GCP    32'h0000000f
`define DCMAC__C0_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_SA_GPP    32'h00000010
`define DCMAC__C0_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_SA_PCP    32'h00000011
`define DCMAC__C0_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_SA_PPP    32'h00000012
`define DCMAC__C0_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_SFD    32'h00000013
`define DCMAC__C0_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_UCAST_GCP    32'h00000014
`define DCMAC__C0_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_UCAST_GPP    32'h00000015
`define DCMAC__C0_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_UCAST_PCP    32'h00000016
`define DCMAC__C0_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C0_CTL_RX_CHECK_UCAST_PPP    32'h00000017
`define DCMAC__C0_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C0_CTL_RX_DATA_RATE    32'h00000018
`define DCMAC__C0_CTL_RX_DATA_RATE_SZ 2

`define DCMAC__C0_CTL_RX_DEGRADE_ACT_THRESH    32'h00000019
`define DCMAC__C0_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C0_CTL_RX_DEGRADE_DEACT_THRESH    32'h0000001a
`define DCMAC__C0_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C0_CTL_RX_DEGRADE_ENABLE    32'h0000001b
`define DCMAC__C0_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C0_CTL_RX_DEGRADE_INTERVAL    32'h0000001c
`define DCMAC__C0_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C0_CTL_RX_DELETE_FCS    32'h0000001d
`define DCMAC__C0_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C0_CTL_RX_ENABLE_GCP    32'h0000001e
`define DCMAC__C0_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C0_CTL_RX_ENABLE_GPP    32'h0000001f
`define DCMAC__C0_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C0_CTL_RX_ENABLE_PCP    32'h00000020
`define DCMAC__C0_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C0_CTL_RX_ENABLE_PPP    32'h00000021
`define DCMAC__C0_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C0_CTL_RX_ETYPE_GCP    32'h00000022
`define DCMAC__C0_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C0_CTL_RX_ETYPE_GPP    32'h00000023
`define DCMAC__C0_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C0_CTL_RX_ETYPE_PCP    32'h00000024
`define DCMAC__C0_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C0_CTL_RX_ETYPE_PPP    32'h00000025
`define DCMAC__C0_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C0_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h00000026
`define DCMAC__C0_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C0_CTL_RX_FEC_BYPASS_CORRECTION    32'h00000027
`define DCMAC__C0_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C0_CTL_RX_FEC_BYPASS_INDICATION    32'h00000028
`define DCMAC__C0_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C0_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h00000029
`define DCMAC__C0_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C0_CTL_RX_FEC_MODE    32'h0000002a
`define DCMAC__C0_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C0_CTL_RX_FEC_TRANSCODE_BYPASS    32'h0000002b
`define DCMAC__C0_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C0_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h0000002c
`define DCMAC__C0_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C0_CTL_RX_FLEXIF_PCS_WIDE_MODE    32'h0000002d
`define DCMAC__C0_CTL_RX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C0_CTL_RX_FLEXIF_SELECT    32'h0000002e
`define DCMAC__C0_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C0_CTL_RX_FORWARD_CONTROL    32'h0000002f
`define DCMAC__C0_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C0_CTL_RX_IGNORE_FCS    32'h00000030
`define DCMAC__C0_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C0_CTL_RX_IGNORE_INRANGE    32'h00000031
`define DCMAC__C0_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C0_CTL_RX_IS_CLAUSE_49    32'h00000032
`define DCMAC__C0_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C0_CTL_RX_MAX_PACKET_LEN    32'h00000033
`define DCMAC__C0_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C0_CTL_RX_OPCODE_GPP    32'h00000034
`define DCMAC__C0_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C0_CTL_RX_OPCODE_MAX_GCP    32'h00000035
`define DCMAC__C0_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C0_CTL_RX_OPCODE_MAX_PCP    32'h00000036
`define DCMAC__C0_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C0_CTL_RX_OPCODE_MIN_GCP    32'h00000037
`define DCMAC__C0_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C0_CTL_RX_OPCODE_MIN_PCP    32'h00000038
`define DCMAC__C0_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C0_CTL_RX_OPCODE_PPP    32'h00000039
`define DCMAC__C0_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C0_CTL_RX_PAUSE_DA_MCAST    32'h0000003a
`define DCMAC__C0_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C0_CTL_RX_PAUSE_DA_UCAST    32'h0000003b
`define DCMAC__C0_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C0_CTL_RX_PAUSE_SA    32'h0000003c
`define DCMAC__C0_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C0_CTL_RX_PMA_LANE_MUX    32'h0000003d
`define DCMAC__C0_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C0_CTL_RX_PROCESS_LFI    32'h0000003e
`define DCMAC__C0_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C0_CTL_RX_PTP_LATENCY_ADJUST    32'h0000003f
`define DCMAC__C0_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C0_CTL_RX_PTP_ST_OFFSET    32'h00000040
`define DCMAC__C0_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C0_CTL_RX_TEST_PATTERN    32'h00000041
`define DCMAC__C0_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C0_CTL_RX_TICK_REG_MODE_SEL    32'h00000042
`define DCMAC__C0_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C0_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000043
`define DCMAC__C0_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C0_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h00000044
`define DCMAC__C0_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C0_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE    32'h00000045
`define DCMAC__C0_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE_SZ 40

`define DCMAC__C0_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000046
`define DCMAC__C0_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C0_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000047
`define DCMAC__C0_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C0_CTL_TX_DATA_RATE    32'h00000048
`define DCMAC__C0_CTL_TX_DATA_RATE_SZ 2

`define DCMAC__C0_CTL_TX_DA_GPP    32'h00000049
`define DCMAC__C0_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C0_CTL_TX_DA_PPP    32'h0000004a
`define DCMAC__C0_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C0_CTL_TX_ETHERTYPE_GPP    32'h0000004b
`define DCMAC__C0_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C0_CTL_TX_ETHERTYPE_PPP    32'h0000004c
`define DCMAC__C0_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C0_CTL_TX_FCS_INS_ENABLE    32'h0000004d
`define DCMAC__C0_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C0_CTL_TX_FEC_FOUR_LANE_PMD    32'h0000004e
`define DCMAC__C0_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C0_CTL_TX_FEC_MODE    32'h0000004f
`define DCMAC__C0_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C0_CTL_TX_FEC_TRANSCODE_BYPASS    32'h00000050
`define DCMAC__C0_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C0_CTL_TX_FLEXIF_AM_MODE    32'h00000051
`define DCMAC__C0_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C0_CTL_TX_FLEXIF_PCS_WIDE_MODE    32'h00000052
`define DCMAC__C0_CTL_TX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C0_CTL_TX_FLEXIF_SELECT    32'h00000053
`define DCMAC__C0_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C0_CTL_TX_IGNORE_FCS    32'h00000054
`define DCMAC__C0_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C0_CTL_TX_IPG_VALUE    32'h00000055
`define DCMAC__C0_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C0_CTL_TX_OPCODE_GPP    32'h00000056
`define DCMAC__C0_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C0_CTL_TX_OPCODE_PPP    32'h00000057
`define DCMAC__C0_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA0    32'h00000058
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA1    32'h00000059
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA2    32'h0000005a
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA3    32'h0000005b
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA4    32'h0000005c
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA5    32'h0000005d
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA6    32'h0000005e
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA7    32'h0000005f
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_QUANTA8    32'h00000060
`define DCMAC__C0_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C0_CTL_TX_PAUSE_REFRESH_TIMER    32'h00000061
`define DCMAC__C0_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C0_CTL_TX_PMA_LANE_MUX    32'h00000062
`define DCMAC__C0_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C0_CTL_TX_PTP_1STEP_ENABLE    32'h00000063
`define DCMAC__C0_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C0_CTL_TX_PTP_LATENCY_ADJUST    32'h00000064
`define DCMAC__C0_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C0_CTL_TX_PTP_SAT_ENABLE    32'h00000065
`define DCMAC__C0_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C0_CTL_TX_PTP_ST_OFFSET    32'h00000066
`define DCMAC__C0_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C0_CTL_TX_SA_GPP    32'h00000067
`define DCMAC__C0_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C0_CTL_TX_SA_PPP    32'h00000068
`define DCMAC__C0_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C0_CTL_TX_SEND_IDLE    32'h00000069
`define DCMAC__C0_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C0_CTL_TX_SEND_LFI    32'h0000006a
`define DCMAC__C0_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C0_CTL_TX_SEND_RFI    32'h0000006b
`define DCMAC__C0_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C0_CTL_TX_TICK_REG_MODE_SEL    32'h0000006c
`define DCMAC__C0_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C0_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h0000006d
`define DCMAC__C0_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C0_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h0000006e
`define DCMAC__C0_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C10_CTL_RX_CHECK_PREAMBLE    32'h0000006f
`define DCMAC__C10_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C10_CTL_RX_CHECK_SFD    32'h00000070
`define DCMAC__C10_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C10_CTL_RX_DELETE_FCS    32'h00000071
`define DCMAC__C10_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C10_CTL_RX_IGNORE_FCS    32'h00000072
`define DCMAC__C10_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C10_CTL_RX_IGNORE_INRANGE    32'h00000073
`define DCMAC__C10_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C10_CTL_RX_IS_CLAUSE_49    32'h00000074
`define DCMAC__C10_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C10_CTL_RX_MAX_PACKET_LEN    32'h00000075
`define DCMAC__C10_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C10_CTL_RX_PROCESS_LFI    32'h00000076
`define DCMAC__C10_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C10_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000077
`define DCMAC__C10_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C10_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000078
`define DCMAC__C10_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C10_CTL_TX_FCS_INS_ENABLE    32'h00000079
`define DCMAC__C10_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C10_CTL_TX_IGNORE_FCS    32'h0000007a
`define DCMAC__C10_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C10_CTL_TX_IPG_VALUE    32'h0000007b
`define DCMAC__C10_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C10_CTL_TX_SEND_IDLE    32'h0000007c
`define DCMAC__C10_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C10_CTL_TX_SEND_LFI    32'h0000007d
`define DCMAC__C10_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C10_CTL_TX_SEND_RFI    32'h0000007e
`define DCMAC__C10_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C11_CTL_RX_CHECK_PREAMBLE    32'h0000007f
`define DCMAC__C11_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C11_CTL_RX_CHECK_SFD    32'h00000080
`define DCMAC__C11_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C11_CTL_RX_DELETE_FCS    32'h00000081
`define DCMAC__C11_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C11_CTL_RX_IGNORE_FCS    32'h00000082
`define DCMAC__C11_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C11_CTL_RX_IGNORE_INRANGE    32'h00000083
`define DCMAC__C11_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C11_CTL_RX_IS_CLAUSE_49    32'h00000084
`define DCMAC__C11_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C11_CTL_RX_MAX_PACKET_LEN    32'h00000085
`define DCMAC__C11_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C11_CTL_RX_PROCESS_LFI    32'h00000086
`define DCMAC__C11_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C11_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000087
`define DCMAC__C11_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C11_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000088
`define DCMAC__C11_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C11_CTL_TX_FCS_INS_ENABLE    32'h00000089
`define DCMAC__C11_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C11_CTL_TX_IGNORE_FCS    32'h0000008a
`define DCMAC__C11_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C11_CTL_TX_IPG_VALUE    32'h0000008b
`define DCMAC__C11_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C11_CTL_TX_SEND_IDLE    32'h0000008c
`define DCMAC__C11_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C11_CTL_TX_SEND_LFI    32'h0000008d
`define DCMAC__C11_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C11_CTL_TX_SEND_RFI    32'h0000008e
`define DCMAC__C11_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C12_CTL_RX_CHECK_PREAMBLE    32'h0000008f
`define DCMAC__C12_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C12_CTL_RX_CHECK_SFD    32'h00000090
`define DCMAC__C12_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C12_CTL_RX_DELETE_FCS    32'h00000091
`define DCMAC__C12_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C12_CTL_RX_IGNORE_FCS    32'h00000092
`define DCMAC__C12_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C12_CTL_RX_IGNORE_INRANGE    32'h00000093
`define DCMAC__C12_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C12_CTL_RX_IS_CLAUSE_49    32'h00000094
`define DCMAC__C12_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C12_CTL_RX_MAX_PACKET_LEN    32'h00000095
`define DCMAC__C12_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C12_CTL_RX_PROCESS_LFI    32'h00000096
`define DCMAC__C12_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C12_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000097
`define DCMAC__C12_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C12_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000098
`define DCMAC__C12_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C12_CTL_TX_FCS_INS_ENABLE    32'h00000099
`define DCMAC__C12_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C12_CTL_TX_IGNORE_FCS    32'h0000009a
`define DCMAC__C12_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C12_CTL_TX_IPG_VALUE    32'h0000009b
`define DCMAC__C12_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C12_CTL_TX_SEND_IDLE    32'h0000009c
`define DCMAC__C12_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C12_CTL_TX_SEND_LFI    32'h0000009d
`define DCMAC__C12_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C12_CTL_TX_SEND_RFI    32'h0000009e
`define DCMAC__C12_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C13_CTL_RX_CHECK_PREAMBLE    32'h0000009f
`define DCMAC__C13_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C13_CTL_RX_CHECK_SFD    32'h000000a0
`define DCMAC__C13_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C13_CTL_RX_DELETE_FCS    32'h000000a1
`define DCMAC__C13_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C13_CTL_RX_IGNORE_FCS    32'h000000a2
`define DCMAC__C13_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C13_CTL_RX_IGNORE_INRANGE    32'h000000a3
`define DCMAC__C13_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C13_CTL_RX_IS_CLAUSE_49    32'h000000a4
`define DCMAC__C13_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C13_CTL_RX_MAX_PACKET_LEN    32'h000000a5
`define DCMAC__C13_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C13_CTL_RX_PROCESS_LFI    32'h000000a6
`define DCMAC__C13_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C13_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000a7
`define DCMAC__C13_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C13_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000a8
`define DCMAC__C13_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C13_CTL_TX_FCS_INS_ENABLE    32'h000000a9
`define DCMAC__C13_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C13_CTL_TX_IGNORE_FCS    32'h000000aa
`define DCMAC__C13_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C13_CTL_TX_IPG_VALUE    32'h000000ab
`define DCMAC__C13_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C13_CTL_TX_SEND_IDLE    32'h000000ac
`define DCMAC__C13_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C13_CTL_TX_SEND_LFI    32'h000000ad
`define DCMAC__C13_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C13_CTL_TX_SEND_RFI    32'h000000ae
`define DCMAC__C13_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C14_CTL_RX_CHECK_PREAMBLE    32'h000000af
`define DCMAC__C14_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C14_CTL_RX_CHECK_SFD    32'h000000b0
`define DCMAC__C14_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C14_CTL_RX_DELETE_FCS    32'h000000b1
`define DCMAC__C14_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C14_CTL_RX_IGNORE_FCS    32'h000000b2
`define DCMAC__C14_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C14_CTL_RX_IGNORE_INRANGE    32'h000000b3
`define DCMAC__C14_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C14_CTL_RX_IS_CLAUSE_49    32'h000000b4
`define DCMAC__C14_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C14_CTL_RX_MAX_PACKET_LEN    32'h000000b5
`define DCMAC__C14_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C14_CTL_RX_PROCESS_LFI    32'h000000b6
`define DCMAC__C14_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C14_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000b7
`define DCMAC__C14_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C14_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000b8
`define DCMAC__C14_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C14_CTL_TX_FCS_INS_ENABLE    32'h000000b9
`define DCMAC__C14_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C14_CTL_TX_IGNORE_FCS    32'h000000ba
`define DCMAC__C14_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C14_CTL_TX_IPG_VALUE    32'h000000bb
`define DCMAC__C14_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C14_CTL_TX_SEND_IDLE    32'h000000bc
`define DCMAC__C14_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C14_CTL_TX_SEND_LFI    32'h000000bd
`define DCMAC__C14_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C14_CTL_TX_SEND_RFI    32'h000000be
`define DCMAC__C14_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C15_CTL_RX_CHECK_PREAMBLE    32'h000000bf
`define DCMAC__C15_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C15_CTL_RX_CHECK_SFD    32'h000000c0
`define DCMAC__C15_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C15_CTL_RX_DELETE_FCS    32'h000000c1
`define DCMAC__C15_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C15_CTL_RX_IGNORE_FCS    32'h000000c2
`define DCMAC__C15_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C15_CTL_RX_IGNORE_INRANGE    32'h000000c3
`define DCMAC__C15_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C15_CTL_RX_IS_CLAUSE_49    32'h000000c4
`define DCMAC__C15_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C15_CTL_RX_MAX_PACKET_LEN    32'h000000c5
`define DCMAC__C15_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C15_CTL_RX_PROCESS_LFI    32'h000000c6
`define DCMAC__C15_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C15_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000c7
`define DCMAC__C15_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C15_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000c8
`define DCMAC__C15_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C15_CTL_TX_FCS_INS_ENABLE    32'h000000c9
`define DCMAC__C15_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C15_CTL_TX_IGNORE_FCS    32'h000000ca
`define DCMAC__C15_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C15_CTL_TX_IPG_VALUE    32'h000000cb
`define DCMAC__C15_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C15_CTL_TX_SEND_IDLE    32'h000000cc
`define DCMAC__C15_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C15_CTL_TX_SEND_LFI    32'h000000cd
`define DCMAC__C15_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C15_CTL_TX_SEND_RFI    32'h000000ce
`define DCMAC__C15_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C16_CTL_RX_CHECK_PREAMBLE    32'h000000cf
`define DCMAC__C16_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C16_CTL_RX_CHECK_SFD    32'h000000d0
`define DCMAC__C16_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C16_CTL_RX_DELETE_FCS    32'h000000d1
`define DCMAC__C16_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C16_CTL_RX_IGNORE_FCS    32'h000000d2
`define DCMAC__C16_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C16_CTL_RX_IGNORE_INRANGE    32'h000000d3
`define DCMAC__C16_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C16_CTL_RX_IS_CLAUSE_49    32'h000000d4
`define DCMAC__C16_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C16_CTL_RX_MAX_PACKET_LEN    32'h000000d5
`define DCMAC__C16_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C16_CTL_RX_PROCESS_LFI    32'h000000d6
`define DCMAC__C16_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C16_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000d7
`define DCMAC__C16_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C16_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000d8
`define DCMAC__C16_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C16_CTL_TX_FCS_INS_ENABLE    32'h000000d9
`define DCMAC__C16_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C16_CTL_TX_IGNORE_FCS    32'h000000da
`define DCMAC__C16_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C16_CTL_TX_IPG_VALUE    32'h000000db
`define DCMAC__C16_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C16_CTL_TX_SEND_IDLE    32'h000000dc
`define DCMAC__C16_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C16_CTL_TX_SEND_LFI    32'h000000dd
`define DCMAC__C16_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C16_CTL_TX_SEND_RFI    32'h000000de
`define DCMAC__C16_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C17_CTL_RX_CHECK_PREAMBLE    32'h000000df
`define DCMAC__C17_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C17_CTL_RX_CHECK_SFD    32'h000000e0
`define DCMAC__C17_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C17_CTL_RX_DELETE_FCS    32'h000000e1
`define DCMAC__C17_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C17_CTL_RX_IGNORE_FCS    32'h000000e2
`define DCMAC__C17_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C17_CTL_RX_IGNORE_INRANGE    32'h000000e3
`define DCMAC__C17_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C17_CTL_RX_IS_CLAUSE_49    32'h000000e4
`define DCMAC__C17_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C17_CTL_RX_MAX_PACKET_LEN    32'h000000e5
`define DCMAC__C17_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C17_CTL_RX_PROCESS_LFI    32'h000000e6
`define DCMAC__C17_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C17_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000e7
`define DCMAC__C17_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C17_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000e8
`define DCMAC__C17_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C17_CTL_TX_FCS_INS_ENABLE    32'h000000e9
`define DCMAC__C17_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C17_CTL_TX_IGNORE_FCS    32'h000000ea
`define DCMAC__C17_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C17_CTL_TX_IPG_VALUE    32'h000000eb
`define DCMAC__C17_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C17_CTL_TX_SEND_IDLE    32'h000000ec
`define DCMAC__C17_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C17_CTL_TX_SEND_LFI    32'h000000ed
`define DCMAC__C17_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C17_CTL_TX_SEND_RFI    32'h000000ee
`define DCMAC__C17_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C18_CTL_RX_CHECK_PREAMBLE    32'h000000ef
`define DCMAC__C18_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C18_CTL_RX_CHECK_SFD    32'h000000f0
`define DCMAC__C18_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C18_CTL_RX_DELETE_FCS    32'h000000f1
`define DCMAC__C18_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C18_CTL_RX_IGNORE_FCS    32'h000000f2
`define DCMAC__C18_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C18_CTL_RX_IGNORE_INRANGE    32'h000000f3
`define DCMAC__C18_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C18_CTL_RX_IS_CLAUSE_49    32'h000000f4
`define DCMAC__C18_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C18_CTL_RX_MAX_PACKET_LEN    32'h000000f5
`define DCMAC__C18_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C18_CTL_RX_PROCESS_LFI    32'h000000f6
`define DCMAC__C18_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C18_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000000f7
`define DCMAC__C18_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C18_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000000f8
`define DCMAC__C18_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C18_CTL_TX_FCS_INS_ENABLE    32'h000000f9
`define DCMAC__C18_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C18_CTL_TX_IGNORE_FCS    32'h000000fa
`define DCMAC__C18_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C18_CTL_TX_IPG_VALUE    32'h000000fb
`define DCMAC__C18_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C18_CTL_TX_SEND_IDLE    32'h000000fc
`define DCMAC__C18_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C18_CTL_TX_SEND_LFI    32'h000000fd
`define DCMAC__C18_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C18_CTL_TX_SEND_RFI    32'h000000fe
`define DCMAC__C18_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C19_CTL_RX_CHECK_PREAMBLE    32'h000000ff
`define DCMAC__C19_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C19_CTL_RX_CHECK_SFD    32'h00000100
`define DCMAC__C19_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C19_CTL_RX_DELETE_FCS    32'h00000101
`define DCMAC__C19_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C19_CTL_RX_IGNORE_FCS    32'h00000102
`define DCMAC__C19_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C19_CTL_RX_IGNORE_INRANGE    32'h00000103
`define DCMAC__C19_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C19_CTL_RX_IS_CLAUSE_49    32'h00000104
`define DCMAC__C19_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C19_CTL_RX_MAX_PACKET_LEN    32'h00000105
`define DCMAC__C19_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C19_CTL_RX_PROCESS_LFI    32'h00000106
`define DCMAC__C19_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C19_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000107
`define DCMAC__C19_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C19_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000108
`define DCMAC__C19_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C19_CTL_TX_FCS_INS_ENABLE    32'h00000109
`define DCMAC__C19_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C19_CTL_TX_IGNORE_FCS    32'h0000010a
`define DCMAC__C19_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C19_CTL_TX_IPG_VALUE    32'h0000010b
`define DCMAC__C19_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C19_CTL_TX_SEND_IDLE    32'h0000010c
`define DCMAC__C19_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C19_CTL_TX_SEND_LFI    32'h0000010d
`define DCMAC__C19_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C19_CTL_TX_SEND_RFI    32'h0000010e
`define DCMAC__C19_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C1_CTL_PCS_RX_TS_EN    32'h0000010f
`define DCMAC__C1_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_ACK    32'h00000110
`define DCMAC__C1_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_ETYPE_GCP    32'h00000111
`define DCMAC__C1_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_ETYPE_GPP    32'h00000112
`define DCMAC__C1_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_ETYPE_PCP    32'h00000113
`define DCMAC__C1_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_ETYPE_PPP    32'h00000114
`define DCMAC__C1_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_MCAST_GCP    32'h00000115
`define DCMAC__C1_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_MCAST_GPP    32'h00000116
`define DCMAC__C1_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_MCAST_PCP    32'h00000117
`define DCMAC__C1_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_MCAST_PPP    32'h00000118
`define DCMAC__C1_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_OPCODE_GCP    32'h00000119
`define DCMAC__C1_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_OPCODE_GPP    32'h0000011a
`define DCMAC__C1_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_OPCODE_PCP    32'h0000011b
`define DCMAC__C1_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_OPCODE_PPP    32'h0000011c
`define DCMAC__C1_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_PREAMBLE    32'h0000011d
`define DCMAC__C1_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_SA_GCP    32'h0000011e
`define DCMAC__C1_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_SA_GPP    32'h0000011f
`define DCMAC__C1_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_SA_PCP    32'h00000120
`define DCMAC__C1_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_SA_PPP    32'h00000121
`define DCMAC__C1_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_SFD    32'h00000122
`define DCMAC__C1_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_UCAST_GCP    32'h00000123
`define DCMAC__C1_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_UCAST_GPP    32'h00000124
`define DCMAC__C1_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_UCAST_PCP    32'h00000125
`define DCMAC__C1_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C1_CTL_RX_CHECK_UCAST_PPP    32'h00000126
`define DCMAC__C1_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C1_CTL_RX_DEGRADE_ACT_THRESH    32'h00000127
`define DCMAC__C1_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C1_CTL_RX_DEGRADE_DEACT_THRESH    32'h00000128
`define DCMAC__C1_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C1_CTL_RX_DEGRADE_ENABLE    32'h00000129
`define DCMAC__C1_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C1_CTL_RX_DEGRADE_INTERVAL    32'h0000012a
`define DCMAC__C1_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C1_CTL_RX_DELETE_FCS    32'h0000012b
`define DCMAC__C1_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C1_CTL_RX_ENABLE_GCP    32'h0000012c
`define DCMAC__C1_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C1_CTL_RX_ENABLE_GPP    32'h0000012d
`define DCMAC__C1_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C1_CTL_RX_ENABLE_PCP    32'h0000012e
`define DCMAC__C1_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C1_CTL_RX_ENABLE_PPP    32'h0000012f
`define DCMAC__C1_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C1_CTL_RX_ETYPE_GCP    32'h00000130
`define DCMAC__C1_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C1_CTL_RX_ETYPE_GPP    32'h00000131
`define DCMAC__C1_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C1_CTL_RX_ETYPE_PCP    32'h00000132
`define DCMAC__C1_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C1_CTL_RX_ETYPE_PPP    32'h00000133
`define DCMAC__C1_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C1_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h00000134
`define DCMAC__C1_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C1_CTL_RX_FEC_BYPASS_CORRECTION    32'h00000135
`define DCMAC__C1_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C1_CTL_RX_FEC_BYPASS_INDICATION    32'h00000136
`define DCMAC__C1_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C1_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h00000137
`define DCMAC__C1_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C1_CTL_RX_FEC_MODE    32'h00000138
`define DCMAC__C1_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C1_CTL_RX_FEC_TRANSCODE_BYPASS    32'h00000139
`define DCMAC__C1_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C1_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h0000013a
`define DCMAC__C1_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C1_CTL_RX_FLEXIF_PCS_WIDE_MODE    32'h0000013b
`define DCMAC__C1_CTL_RX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C1_CTL_RX_FLEXIF_SELECT    32'h0000013c
`define DCMAC__C1_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C1_CTL_RX_FORWARD_CONTROL    32'h0000013d
`define DCMAC__C1_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C1_CTL_RX_IGNORE_FCS    32'h0000013e
`define DCMAC__C1_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C1_CTL_RX_IGNORE_INRANGE    32'h0000013f
`define DCMAC__C1_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C1_CTL_RX_IS_CLAUSE_49    32'h00000140
`define DCMAC__C1_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C1_CTL_RX_MAX_PACKET_LEN    32'h00000141
`define DCMAC__C1_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C1_CTL_RX_OPCODE_GPP    32'h00000142
`define DCMAC__C1_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C1_CTL_RX_OPCODE_MAX_GCP    32'h00000143
`define DCMAC__C1_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C1_CTL_RX_OPCODE_MAX_PCP    32'h00000144
`define DCMAC__C1_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C1_CTL_RX_OPCODE_MIN_GCP    32'h00000145
`define DCMAC__C1_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C1_CTL_RX_OPCODE_MIN_PCP    32'h00000146
`define DCMAC__C1_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C1_CTL_RX_OPCODE_PPP    32'h00000147
`define DCMAC__C1_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C1_CTL_RX_PAUSE_DA_MCAST    32'h00000148
`define DCMAC__C1_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C1_CTL_RX_PAUSE_DA_UCAST    32'h00000149
`define DCMAC__C1_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C1_CTL_RX_PAUSE_SA    32'h0000014a
`define DCMAC__C1_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C1_CTL_RX_PMA_LANE_MUX    32'h0000014b
`define DCMAC__C1_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C1_CTL_RX_PROCESS_LFI    32'h0000014c
`define DCMAC__C1_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C1_CTL_RX_PTP_LATENCY_ADJUST    32'h0000014d
`define DCMAC__C1_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C1_CTL_RX_PTP_ST_OFFSET    32'h0000014e
`define DCMAC__C1_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C1_CTL_RX_TEST_PATTERN    32'h0000014f
`define DCMAC__C1_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C1_CTL_RX_TICK_REG_MODE_SEL    32'h00000150
`define DCMAC__C1_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C1_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000151
`define DCMAC__C1_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C1_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h00000152
`define DCMAC__C1_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C1_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000153
`define DCMAC__C1_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C1_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000154
`define DCMAC__C1_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C1_CTL_TX_DA_GPP    32'h00000155
`define DCMAC__C1_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C1_CTL_TX_DA_PPP    32'h00000156
`define DCMAC__C1_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C1_CTL_TX_ETHERTYPE_GPP    32'h00000157
`define DCMAC__C1_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C1_CTL_TX_ETHERTYPE_PPP    32'h00000158
`define DCMAC__C1_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C1_CTL_TX_FCS_INS_ENABLE    32'h00000159
`define DCMAC__C1_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C1_CTL_TX_FEC_FOUR_LANE_PMD    32'h0000015a
`define DCMAC__C1_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C1_CTL_TX_FEC_MODE    32'h0000015b
`define DCMAC__C1_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C1_CTL_TX_FEC_TRANSCODE_BYPASS    32'h0000015c
`define DCMAC__C1_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C1_CTL_TX_FLEXIF_AM_MODE    32'h0000015d
`define DCMAC__C1_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C1_CTL_TX_FLEXIF_PCS_WIDE_MODE    32'h0000015e
`define DCMAC__C1_CTL_TX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C1_CTL_TX_FLEXIF_SELECT    32'h0000015f
`define DCMAC__C1_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C1_CTL_TX_IGNORE_FCS    32'h00000160
`define DCMAC__C1_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C1_CTL_TX_IPG_VALUE    32'h00000161
`define DCMAC__C1_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C1_CTL_TX_OPCODE_GPP    32'h00000162
`define DCMAC__C1_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C1_CTL_TX_OPCODE_PPP    32'h00000163
`define DCMAC__C1_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA0    32'h00000164
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA1    32'h00000165
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA2    32'h00000166
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA3    32'h00000167
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA4    32'h00000168
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA5    32'h00000169
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA6    32'h0000016a
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA7    32'h0000016b
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_QUANTA8    32'h0000016c
`define DCMAC__C1_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C1_CTL_TX_PAUSE_REFRESH_TIMER    32'h0000016d
`define DCMAC__C1_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C1_CTL_TX_PMA_LANE_MUX    32'h0000016e
`define DCMAC__C1_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C1_CTL_TX_PTP_1STEP_ENABLE    32'h0000016f
`define DCMAC__C1_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C1_CTL_TX_PTP_LATENCY_ADJUST    32'h00000170
`define DCMAC__C1_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C1_CTL_TX_PTP_SAT_ENABLE    32'h00000171
`define DCMAC__C1_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C1_CTL_TX_PTP_ST_OFFSET    32'h00000172
`define DCMAC__C1_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C1_CTL_TX_SA_GPP    32'h00000173
`define DCMAC__C1_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C1_CTL_TX_SA_PPP    32'h00000174
`define DCMAC__C1_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C1_CTL_TX_SEND_IDLE    32'h00000175
`define DCMAC__C1_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C1_CTL_TX_SEND_LFI    32'h00000176
`define DCMAC__C1_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C1_CTL_TX_SEND_RFI    32'h00000177
`define DCMAC__C1_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C1_CTL_TX_TICK_REG_MODE_SEL    32'h00000178
`define DCMAC__C1_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C1_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000179
`define DCMAC__C1_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C1_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h0000017a
`define DCMAC__C1_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C20_CTL_RX_CHECK_PREAMBLE    32'h0000017b
`define DCMAC__C20_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C20_CTL_RX_CHECK_SFD    32'h0000017c
`define DCMAC__C20_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C20_CTL_RX_DELETE_FCS    32'h0000017d
`define DCMAC__C20_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C20_CTL_RX_IGNORE_FCS    32'h0000017e
`define DCMAC__C20_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C20_CTL_RX_IGNORE_INRANGE    32'h0000017f
`define DCMAC__C20_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C20_CTL_RX_IS_CLAUSE_49    32'h00000180
`define DCMAC__C20_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C20_CTL_RX_MAX_PACKET_LEN    32'h00000181
`define DCMAC__C20_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C20_CTL_RX_PROCESS_LFI    32'h00000182
`define DCMAC__C20_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C20_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000183
`define DCMAC__C20_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C20_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000184
`define DCMAC__C20_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C20_CTL_TX_FCS_INS_ENABLE    32'h00000185
`define DCMAC__C20_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C20_CTL_TX_IGNORE_FCS    32'h00000186
`define DCMAC__C20_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C20_CTL_TX_IPG_VALUE    32'h00000187
`define DCMAC__C20_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C20_CTL_TX_SEND_IDLE    32'h00000188
`define DCMAC__C20_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C20_CTL_TX_SEND_LFI    32'h00000189
`define DCMAC__C20_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C20_CTL_TX_SEND_RFI    32'h0000018a
`define DCMAC__C20_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C21_CTL_RX_CHECK_PREAMBLE    32'h0000018b
`define DCMAC__C21_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C21_CTL_RX_CHECK_SFD    32'h0000018c
`define DCMAC__C21_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C21_CTL_RX_DELETE_FCS    32'h0000018d
`define DCMAC__C21_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C21_CTL_RX_IGNORE_FCS    32'h0000018e
`define DCMAC__C21_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C21_CTL_RX_IGNORE_INRANGE    32'h0000018f
`define DCMAC__C21_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C21_CTL_RX_IS_CLAUSE_49    32'h00000190
`define DCMAC__C21_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C21_CTL_RX_MAX_PACKET_LEN    32'h00000191
`define DCMAC__C21_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C21_CTL_RX_PROCESS_LFI    32'h00000192
`define DCMAC__C21_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C21_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000193
`define DCMAC__C21_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C21_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000194
`define DCMAC__C21_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C21_CTL_TX_FCS_INS_ENABLE    32'h00000195
`define DCMAC__C21_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C21_CTL_TX_IGNORE_FCS    32'h00000196
`define DCMAC__C21_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C21_CTL_TX_IPG_VALUE    32'h00000197
`define DCMAC__C21_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C21_CTL_TX_SEND_IDLE    32'h00000198
`define DCMAC__C21_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C21_CTL_TX_SEND_LFI    32'h00000199
`define DCMAC__C21_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C21_CTL_TX_SEND_RFI    32'h0000019a
`define DCMAC__C21_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C22_CTL_RX_CHECK_PREAMBLE    32'h0000019b
`define DCMAC__C22_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C22_CTL_RX_CHECK_SFD    32'h0000019c
`define DCMAC__C22_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C22_CTL_RX_DELETE_FCS    32'h0000019d
`define DCMAC__C22_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C22_CTL_RX_IGNORE_FCS    32'h0000019e
`define DCMAC__C22_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C22_CTL_RX_IGNORE_INRANGE    32'h0000019f
`define DCMAC__C22_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C22_CTL_RX_IS_CLAUSE_49    32'h000001a0
`define DCMAC__C22_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C22_CTL_RX_MAX_PACKET_LEN    32'h000001a1
`define DCMAC__C22_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C22_CTL_RX_PROCESS_LFI    32'h000001a2
`define DCMAC__C22_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C22_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001a3
`define DCMAC__C22_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C22_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001a4
`define DCMAC__C22_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C22_CTL_TX_FCS_INS_ENABLE    32'h000001a5
`define DCMAC__C22_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C22_CTL_TX_IGNORE_FCS    32'h000001a6
`define DCMAC__C22_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C22_CTL_TX_IPG_VALUE    32'h000001a7
`define DCMAC__C22_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C22_CTL_TX_SEND_IDLE    32'h000001a8
`define DCMAC__C22_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C22_CTL_TX_SEND_LFI    32'h000001a9
`define DCMAC__C22_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C22_CTL_TX_SEND_RFI    32'h000001aa
`define DCMAC__C22_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C23_CTL_RX_CHECK_PREAMBLE    32'h000001ab
`define DCMAC__C23_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C23_CTL_RX_CHECK_SFD    32'h000001ac
`define DCMAC__C23_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C23_CTL_RX_DELETE_FCS    32'h000001ad
`define DCMAC__C23_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C23_CTL_RX_IGNORE_FCS    32'h000001ae
`define DCMAC__C23_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C23_CTL_RX_IGNORE_INRANGE    32'h000001af
`define DCMAC__C23_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C23_CTL_RX_IS_CLAUSE_49    32'h000001b0
`define DCMAC__C23_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C23_CTL_RX_MAX_PACKET_LEN    32'h000001b1
`define DCMAC__C23_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C23_CTL_RX_PROCESS_LFI    32'h000001b2
`define DCMAC__C23_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C23_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001b3
`define DCMAC__C23_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C23_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001b4
`define DCMAC__C23_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C23_CTL_TX_FCS_INS_ENABLE    32'h000001b5
`define DCMAC__C23_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C23_CTL_TX_IGNORE_FCS    32'h000001b6
`define DCMAC__C23_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C23_CTL_TX_IPG_VALUE    32'h000001b7
`define DCMAC__C23_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C23_CTL_TX_SEND_IDLE    32'h000001b8
`define DCMAC__C23_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C23_CTL_TX_SEND_LFI    32'h000001b9
`define DCMAC__C23_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C23_CTL_TX_SEND_RFI    32'h000001ba
`define DCMAC__C23_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C24_CTL_RX_CHECK_PREAMBLE    32'h000001bb
`define DCMAC__C24_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C24_CTL_RX_CHECK_SFD    32'h000001bc
`define DCMAC__C24_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C24_CTL_RX_DELETE_FCS    32'h000001bd
`define DCMAC__C24_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C24_CTL_RX_IGNORE_FCS    32'h000001be
`define DCMAC__C24_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C24_CTL_RX_IGNORE_INRANGE    32'h000001bf
`define DCMAC__C24_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C24_CTL_RX_IS_CLAUSE_49    32'h000001c0
`define DCMAC__C24_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C24_CTL_RX_MAX_PACKET_LEN    32'h000001c1
`define DCMAC__C24_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C24_CTL_RX_PROCESS_LFI    32'h000001c2
`define DCMAC__C24_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C24_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001c3
`define DCMAC__C24_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C24_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001c4
`define DCMAC__C24_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C24_CTL_TX_FCS_INS_ENABLE    32'h000001c5
`define DCMAC__C24_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C24_CTL_TX_IGNORE_FCS    32'h000001c6
`define DCMAC__C24_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C24_CTL_TX_IPG_VALUE    32'h000001c7
`define DCMAC__C24_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C24_CTL_TX_SEND_IDLE    32'h000001c8
`define DCMAC__C24_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C24_CTL_TX_SEND_LFI    32'h000001c9
`define DCMAC__C24_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C24_CTL_TX_SEND_RFI    32'h000001ca
`define DCMAC__C24_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C25_CTL_RX_CHECK_PREAMBLE    32'h000001cb
`define DCMAC__C25_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C25_CTL_RX_CHECK_SFD    32'h000001cc
`define DCMAC__C25_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C25_CTL_RX_DELETE_FCS    32'h000001cd
`define DCMAC__C25_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C25_CTL_RX_IGNORE_FCS    32'h000001ce
`define DCMAC__C25_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C25_CTL_RX_IGNORE_INRANGE    32'h000001cf
`define DCMAC__C25_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C25_CTL_RX_IS_CLAUSE_49    32'h000001d0
`define DCMAC__C25_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C25_CTL_RX_MAX_PACKET_LEN    32'h000001d1
`define DCMAC__C25_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C25_CTL_RX_PROCESS_LFI    32'h000001d2
`define DCMAC__C25_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C25_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001d3
`define DCMAC__C25_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C25_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001d4
`define DCMAC__C25_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C25_CTL_TX_FCS_INS_ENABLE    32'h000001d5
`define DCMAC__C25_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C25_CTL_TX_IGNORE_FCS    32'h000001d6
`define DCMAC__C25_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C25_CTL_TX_IPG_VALUE    32'h000001d7
`define DCMAC__C25_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C25_CTL_TX_SEND_IDLE    32'h000001d8
`define DCMAC__C25_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C25_CTL_TX_SEND_LFI    32'h000001d9
`define DCMAC__C25_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C25_CTL_TX_SEND_RFI    32'h000001da
`define DCMAC__C25_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C26_CTL_RX_CHECK_PREAMBLE    32'h000001db
`define DCMAC__C26_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C26_CTL_RX_CHECK_SFD    32'h000001dc
`define DCMAC__C26_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C26_CTL_RX_DELETE_FCS    32'h000001dd
`define DCMAC__C26_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C26_CTL_RX_IGNORE_FCS    32'h000001de
`define DCMAC__C26_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C26_CTL_RX_IGNORE_INRANGE    32'h000001df
`define DCMAC__C26_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C26_CTL_RX_IS_CLAUSE_49    32'h000001e0
`define DCMAC__C26_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C26_CTL_RX_MAX_PACKET_LEN    32'h000001e1
`define DCMAC__C26_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C26_CTL_RX_PROCESS_LFI    32'h000001e2
`define DCMAC__C26_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C26_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001e3
`define DCMAC__C26_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C26_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001e4
`define DCMAC__C26_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C26_CTL_TX_FCS_INS_ENABLE    32'h000001e5
`define DCMAC__C26_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C26_CTL_TX_IGNORE_FCS    32'h000001e6
`define DCMAC__C26_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C26_CTL_TX_IPG_VALUE    32'h000001e7
`define DCMAC__C26_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C26_CTL_TX_SEND_IDLE    32'h000001e8
`define DCMAC__C26_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C26_CTL_TX_SEND_LFI    32'h000001e9
`define DCMAC__C26_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C26_CTL_TX_SEND_RFI    32'h000001ea
`define DCMAC__C26_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C27_CTL_RX_CHECK_PREAMBLE    32'h000001eb
`define DCMAC__C27_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C27_CTL_RX_CHECK_SFD    32'h000001ec
`define DCMAC__C27_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C27_CTL_RX_DELETE_FCS    32'h000001ed
`define DCMAC__C27_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C27_CTL_RX_IGNORE_FCS    32'h000001ee
`define DCMAC__C27_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C27_CTL_RX_IGNORE_INRANGE    32'h000001ef
`define DCMAC__C27_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C27_CTL_RX_IS_CLAUSE_49    32'h000001f0
`define DCMAC__C27_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C27_CTL_RX_MAX_PACKET_LEN    32'h000001f1
`define DCMAC__C27_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C27_CTL_RX_PROCESS_LFI    32'h000001f2
`define DCMAC__C27_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C27_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000001f3
`define DCMAC__C27_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C27_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000001f4
`define DCMAC__C27_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C27_CTL_TX_FCS_INS_ENABLE    32'h000001f5
`define DCMAC__C27_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C27_CTL_TX_IGNORE_FCS    32'h000001f6
`define DCMAC__C27_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C27_CTL_TX_IPG_VALUE    32'h000001f7
`define DCMAC__C27_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C27_CTL_TX_SEND_IDLE    32'h000001f8
`define DCMAC__C27_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C27_CTL_TX_SEND_LFI    32'h000001f9
`define DCMAC__C27_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C27_CTL_TX_SEND_RFI    32'h000001fa
`define DCMAC__C27_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C28_CTL_RX_CHECK_PREAMBLE    32'h000001fb
`define DCMAC__C28_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C28_CTL_RX_CHECK_SFD    32'h000001fc
`define DCMAC__C28_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C28_CTL_RX_DELETE_FCS    32'h000001fd
`define DCMAC__C28_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C28_CTL_RX_IGNORE_FCS    32'h000001fe
`define DCMAC__C28_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C28_CTL_RX_IGNORE_INRANGE    32'h000001ff
`define DCMAC__C28_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C28_CTL_RX_IS_CLAUSE_49    32'h00000200
`define DCMAC__C28_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C28_CTL_RX_MAX_PACKET_LEN    32'h00000201
`define DCMAC__C28_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C28_CTL_RX_PROCESS_LFI    32'h00000202
`define DCMAC__C28_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C28_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000203
`define DCMAC__C28_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C28_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000204
`define DCMAC__C28_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C28_CTL_TX_FCS_INS_ENABLE    32'h00000205
`define DCMAC__C28_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C28_CTL_TX_IGNORE_FCS    32'h00000206
`define DCMAC__C28_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C28_CTL_TX_IPG_VALUE    32'h00000207
`define DCMAC__C28_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C28_CTL_TX_SEND_IDLE    32'h00000208
`define DCMAC__C28_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C28_CTL_TX_SEND_LFI    32'h00000209
`define DCMAC__C28_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C28_CTL_TX_SEND_RFI    32'h0000020a
`define DCMAC__C28_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C29_CTL_RX_CHECK_PREAMBLE    32'h0000020b
`define DCMAC__C29_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C29_CTL_RX_CHECK_SFD    32'h0000020c
`define DCMAC__C29_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C29_CTL_RX_DELETE_FCS    32'h0000020d
`define DCMAC__C29_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C29_CTL_RX_IGNORE_FCS    32'h0000020e
`define DCMAC__C29_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C29_CTL_RX_IGNORE_INRANGE    32'h0000020f
`define DCMAC__C29_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C29_CTL_RX_IS_CLAUSE_49    32'h00000210
`define DCMAC__C29_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C29_CTL_RX_MAX_PACKET_LEN    32'h00000211
`define DCMAC__C29_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C29_CTL_RX_PROCESS_LFI    32'h00000212
`define DCMAC__C29_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C29_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000213
`define DCMAC__C29_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C29_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000214
`define DCMAC__C29_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C29_CTL_TX_FCS_INS_ENABLE    32'h00000215
`define DCMAC__C29_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C29_CTL_TX_IGNORE_FCS    32'h00000216
`define DCMAC__C29_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C29_CTL_TX_IPG_VALUE    32'h00000217
`define DCMAC__C29_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C29_CTL_TX_SEND_IDLE    32'h00000218
`define DCMAC__C29_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C29_CTL_TX_SEND_LFI    32'h00000219
`define DCMAC__C29_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C29_CTL_TX_SEND_RFI    32'h0000021a
`define DCMAC__C29_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C2_CTL_PCS_RX_TS_EN    32'h0000021b
`define DCMAC__C2_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_ACK    32'h0000021c
`define DCMAC__C2_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_ETYPE_GCP    32'h0000021d
`define DCMAC__C2_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_ETYPE_GPP    32'h0000021e
`define DCMAC__C2_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_ETYPE_PCP    32'h0000021f
`define DCMAC__C2_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_ETYPE_PPP    32'h00000220
`define DCMAC__C2_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_MCAST_GCP    32'h00000221
`define DCMAC__C2_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_MCAST_GPP    32'h00000222
`define DCMAC__C2_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_MCAST_PCP    32'h00000223
`define DCMAC__C2_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_MCAST_PPP    32'h00000224
`define DCMAC__C2_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_OPCODE_GCP    32'h00000225
`define DCMAC__C2_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_OPCODE_GPP    32'h00000226
`define DCMAC__C2_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_OPCODE_PCP    32'h00000227
`define DCMAC__C2_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_OPCODE_PPP    32'h00000228
`define DCMAC__C2_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_PREAMBLE    32'h00000229
`define DCMAC__C2_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_SA_GCP    32'h0000022a
`define DCMAC__C2_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_SA_GPP    32'h0000022b
`define DCMAC__C2_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_SA_PCP    32'h0000022c
`define DCMAC__C2_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_SA_PPP    32'h0000022d
`define DCMAC__C2_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_SFD    32'h0000022e
`define DCMAC__C2_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_UCAST_GCP    32'h0000022f
`define DCMAC__C2_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_UCAST_GPP    32'h00000230
`define DCMAC__C2_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_UCAST_PCP    32'h00000231
`define DCMAC__C2_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C2_CTL_RX_CHECK_UCAST_PPP    32'h00000232
`define DCMAC__C2_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C2_CTL_RX_DATA_RATE    32'h00000233
`define DCMAC__C2_CTL_RX_DATA_RATE_SZ 1

`define DCMAC__C2_CTL_RX_DEGRADE_ACT_THRESH    32'h00000234
`define DCMAC__C2_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C2_CTL_RX_DEGRADE_DEACT_THRESH    32'h00000235
`define DCMAC__C2_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C2_CTL_RX_DEGRADE_ENABLE    32'h00000236
`define DCMAC__C2_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C2_CTL_RX_DEGRADE_INTERVAL    32'h00000237
`define DCMAC__C2_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C2_CTL_RX_DELETE_FCS    32'h00000238
`define DCMAC__C2_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C2_CTL_RX_ENABLE_GCP    32'h00000239
`define DCMAC__C2_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C2_CTL_RX_ENABLE_GPP    32'h0000023a
`define DCMAC__C2_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C2_CTL_RX_ENABLE_PCP    32'h0000023b
`define DCMAC__C2_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C2_CTL_RX_ENABLE_PPP    32'h0000023c
`define DCMAC__C2_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C2_CTL_RX_ETYPE_GCP    32'h0000023d
`define DCMAC__C2_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C2_CTL_RX_ETYPE_GPP    32'h0000023e
`define DCMAC__C2_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C2_CTL_RX_ETYPE_PCP    32'h0000023f
`define DCMAC__C2_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C2_CTL_RX_ETYPE_PPP    32'h00000240
`define DCMAC__C2_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C2_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h00000241
`define DCMAC__C2_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C2_CTL_RX_FEC_BYPASS_CORRECTION    32'h00000242
`define DCMAC__C2_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C2_CTL_RX_FEC_BYPASS_INDICATION    32'h00000243
`define DCMAC__C2_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C2_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h00000244
`define DCMAC__C2_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C2_CTL_RX_FEC_MODE    32'h00000245
`define DCMAC__C2_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C2_CTL_RX_FEC_TRANSCODE_BYPASS    32'h00000246
`define DCMAC__C2_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C2_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h00000247
`define DCMAC__C2_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C2_CTL_RX_FLEXIF_PCS_WIDE_MODE    32'h00000248
`define DCMAC__C2_CTL_RX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C2_CTL_RX_FLEXIF_SELECT    32'h00000249
`define DCMAC__C2_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C2_CTL_RX_FORWARD_CONTROL    32'h0000024a
`define DCMAC__C2_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C2_CTL_RX_IGNORE_FCS    32'h0000024b
`define DCMAC__C2_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C2_CTL_RX_IGNORE_INRANGE    32'h0000024c
`define DCMAC__C2_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C2_CTL_RX_IS_CLAUSE_49    32'h0000024d
`define DCMAC__C2_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C2_CTL_RX_MAX_PACKET_LEN    32'h0000024e
`define DCMAC__C2_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C2_CTL_RX_OPCODE_GPP    32'h0000024f
`define DCMAC__C2_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C2_CTL_RX_OPCODE_MAX_GCP    32'h00000250
`define DCMAC__C2_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C2_CTL_RX_OPCODE_MAX_PCP    32'h00000251
`define DCMAC__C2_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C2_CTL_RX_OPCODE_MIN_GCP    32'h00000252
`define DCMAC__C2_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C2_CTL_RX_OPCODE_MIN_PCP    32'h00000253
`define DCMAC__C2_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C2_CTL_RX_OPCODE_PPP    32'h00000254
`define DCMAC__C2_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C2_CTL_RX_PAUSE_DA_MCAST    32'h00000255
`define DCMAC__C2_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C2_CTL_RX_PAUSE_DA_UCAST    32'h00000256
`define DCMAC__C2_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C2_CTL_RX_PAUSE_SA    32'h00000257
`define DCMAC__C2_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C2_CTL_RX_PMA_LANE_MUX    32'h00000258
`define DCMAC__C2_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C2_CTL_RX_PROCESS_LFI    32'h00000259
`define DCMAC__C2_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C2_CTL_RX_PTP_LATENCY_ADJUST    32'h0000025a
`define DCMAC__C2_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C2_CTL_RX_PTP_ST_OFFSET    32'h0000025b
`define DCMAC__C2_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C2_CTL_RX_TEST_PATTERN    32'h0000025c
`define DCMAC__C2_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C2_CTL_RX_TICK_REG_MODE_SEL    32'h0000025d
`define DCMAC__C2_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C2_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h0000025e
`define DCMAC__C2_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C2_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h0000025f
`define DCMAC__C2_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C2_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE    32'h00000260
`define DCMAC__C2_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE_SZ 40

`define DCMAC__C2_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000261
`define DCMAC__C2_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C2_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000262
`define DCMAC__C2_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C2_CTL_TX_DATA_RATE    32'h00000263
`define DCMAC__C2_CTL_TX_DATA_RATE_SZ 1

`define DCMAC__C2_CTL_TX_DA_GPP    32'h00000264
`define DCMAC__C2_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C2_CTL_TX_DA_PPP    32'h00000265
`define DCMAC__C2_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C2_CTL_TX_ETHERTYPE_GPP    32'h00000266
`define DCMAC__C2_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C2_CTL_TX_ETHERTYPE_PPP    32'h00000267
`define DCMAC__C2_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C2_CTL_TX_FCS_INS_ENABLE    32'h00000268
`define DCMAC__C2_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C2_CTL_TX_FEC_FOUR_LANE_PMD    32'h00000269
`define DCMAC__C2_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C2_CTL_TX_FEC_MODE    32'h0000026a
`define DCMAC__C2_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C2_CTL_TX_FEC_TRANSCODE_BYPASS    32'h0000026b
`define DCMAC__C2_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C2_CTL_TX_FLEXIF_AM_MODE    32'h0000026c
`define DCMAC__C2_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C2_CTL_TX_FLEXIF_PCS_WIDE_MODE    32'h0000026d
`define DCMAC__C2_CTL_TX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C2_CTL_TX_FLEXIF_SELECT    32'h0000026e
`define DCMAC__C2_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C2_CTL_TX_IGNORE_FCS    32'h0000026f
`define DCMAC__C2_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C2_CTL_TX_IPG_VALUE    32'h00000270
`define DCMAC__C2_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C2_CTL_TX_OPCODE_GPP    32'h00000271
`define DCMAC__C2_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C2_CTL_TX_OPCODE_PPP    32'h00000272
`define DCMAC__C2_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA0    32'h00000273
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA1    32'h00000274
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA2    32'h00000275
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA3    32'h00000276
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA4    32'h00000277
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA5    32'h00000278
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA6    32'h00000279
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA7    32'h0000027a
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_QUANTA8    32'h0000027b
`define DCMAC__C2_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C2_CTL_TX_PAUSE_REFRESH_TIMER    32'h0000027c
`define DCMAC__C2_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C2_CTL_TX_PMA_LANE_MUX    32'h0000027d
`define DCMAC__C2_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C2_CTL_TX_PTP_1STEP_ENABLE    32'h0000027e
`define DCMAC__C2_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C2_CTL_TX_PTP_LATENCY_ADJUST    32'h0000027f
`define DCMAC__C2_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C2_CTL_TX_PTP_SAT_ENABLE    32'h00000280
`define DCMAC__C2_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C2_CTL_TX_PTP_ST_OFFSET    32'h00000281
`define DCMAC__C2_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C2_CTL_TX_SA_GPP    32'h00000282
`define DCMAC__C2_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C2_CTL_TX_SA_PPP    32'h00000283
`define DCMAC__C2_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C2_CTL_TX_SEND_IDLE    32'h00000284
`define DCMAC__C2_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C2_CTL_TX_SEND_LFI    32'h00000285
`define DCMAC__C2_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C2_CTL_TX_SEND_RFI    32'h00000286
`define DCMAC__C2_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C2_CTL_TX_TICK_REG_MODE_SEL    32'h00000287
`define DCMAC__C2_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C2_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000288
`define DCMAC__C2_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C2_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h00000289
`define DCMAC__C2_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C30_CTL_RX_CHECK_PREAMBLE    32'h0000028a
`define DCMAC__C30_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C30_CTL_RX_CHECK_SFD    32'h0000028b
`define DCMAC__C30_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C30_CTL_RX_DELETE_FCS    32'h0000028c
`define DCMAC__C30_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C30_CTL_RX_IGNORE_FCS    32'h0000028d
`define DCMAC__C30_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C30_CTL_RX_IGNORE_INRANGE    32'h0000028e
`define DCMAC__C30_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C30_CTL_RX_IS_CLAUSE_49    32'h0000028f
`define DCMAC__C30_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C30_CTL_RX_MAX_PACKET_LEN    32'h00000290
`define DCMAC__C30_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C30_CTL_RX_PROCESS_LFI    32'h00000291
`define DCMAC__C30_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C30_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000292
`define DCMAC__C30_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C30_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000293
`define DCMAC__C30_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C30_CTL_TX_FCS_INS_ENABLE    32'h00000294
`define DCMAC__C30_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C30_CTL_TX_IGNORE_FCS    32'h00000295
`define DCMAC__C30_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C30_CTL_TX_IPG_VALUE    32'h00000296
`define DCMAC__C30_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C30_CTL_TX_SEND_IDLE    32'h00000297
`define DCMAC__C30_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C30_CTL_TX_SEND_LFI    32'h00000298
`define DCMAC__C30_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C30_CTL_TX_SEND_RFI    32'h00000299
`define DCMAC__C30_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C31_CTL_RX_CHECK_PREAMBLE    32'h0000029a
`define DCMAC__C31_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C31_CTL_RX_CHECK_SFD    32'h0000029b
`define DCMAC__C31_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C31_CTL_RX_DELETE_FCS    32'h0000029c
`define DCMAC__C31_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C31_CTL_RX_IGNORE_FCS    32'h0000029d
`define DCMAC__C31_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C31_CTL_RX_IGNORE_INRANGE    32'h0000029e
`define DCMAC__C31_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C31_CTL_RX_IS_CLAUSE_49    32'h0000029f
`define DCMAC__C31_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C31_CTL_RX_MAX_PACKET_LEN    32'h000002a0
`define DCMAC__C31_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C31_CTL_RX_PROCESS_LFI    32'h000002a1
`define DCMAC__C31_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C31_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002a2
`define DCMAC__C31_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C31_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002a3
`define DCMAC__C31_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C31_CTL_TX_FCS_INS_ENABLE    32'h000002a4
`define DCMAC__C31_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C31_CTL_TX_IGNORE_FCS    32'h000002a5
`define DCMAC__C31_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C31_CTL_TX_IPG_VALUE    32'h000002a6
`define DCMAC__C31_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C31_CTL_TX_SEND_IDLE    32'h000002a7
`define DCMAC__C31_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C31_CTL_TX_SEND_LFI    32'h000002a8
`define DCMAC__C31_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C31_CTL_TX_SEND_RFI    32'h000002a9
`define DCMAC__C31_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C32_CTL_RX_CHECK_PREAMBLE    32'h000002aa
`define DCMAC__C32_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C32_CTL_RX_CHECK_SFD    32'h000002ab
`define DCMAC__C32_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C32_CTL_RX_DELETE_FCS    32'h000002ac
`define DCMAC__C32_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C32_CTL_RX_IGNORE_FCS    32'h000002ad
`define DCMAC__C32_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C32_CTL_RX_IGNORE_INRANGE    32'h000002ae
`define DCMAC__C32_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C32_CTL_RX_IS_CLAUSE_49    32'h000002af
`define DCMAC__C32_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C32_CTL_RX_MAX_PACKET_LEN    32'h000002b0
`define DCMAC__C32_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C32_CTL_RX_PROCESS_LFI    32'h000002b1
`define DCMAC__C32_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C32_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002b2
`define DCMAC__C32_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C32_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002b3
`define DCMAC__C32_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C32_CTL_TX_FCS_INS_ENABLE    32'h000002b4
`define DCMAC__C32_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C32_CTL_TX_IGNORE_FCS    32'h000002b5
`define DCMAC__C32_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C32_CTL_TX_IPG_VALUE    32'h000002b6
`define DCMAC__C32_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C32_CTL_TX_SEND_IDLE    32'h000002b7
`define DCMAC__C32_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C32_CTL_TX_SEND_LFI    32'h000002b8
`define DCMAC__C32_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C32_CTL_TX_SEND_RFI    32'h000002b9
`define DCMAC__C32_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C33_CTL_RX_CHECK_PREAMBLE    32'h000002ba
`define DCMAC__C33_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C33_CTL_RX_CHECK_SFD    32'h000002bb
`define DCMAC__C33_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C33_CTL_RX_DELETE_FCS    32'h000002bc
`define DCMAC__C33_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C33_CTL_RX_IGNORE_FCS    32'h000002bd
`define DCMAC__C33_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C33_CTL_RX_IGNORE_INRANGE    32'h000002be
`define DCMAC__C33_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C33_CTL_RX_IS_CLAUSE_49    32'h000002bf
`define DCMAC__C33_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C33_CTL_RX_MAX_PACKET_LEN    32'h000002c0
`define DCMAC__C33_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C33_CTL_RX_PROCESS_LFI    32'h000002c1
`define DCMAC__C33_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C33_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002c2
`define DCMAC__C33_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C33_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002c3
`define DCMAC__C33_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C33_CTL_TX_FCS_INS_ENABLE    32'h000002c4
`define DCMAC__C33_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C33_CTL_TX_IGNORE_FCS    32'h000002c5
`define DCMAC__C33_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C33_CTL_TX_IPG_VALUE    32'h000002c6
`define DCMAC__C33_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C33_CTL_TX_SEND_IDLE    32'h000002c7
`define DCMAC__C33_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C33_CTL_TX_SEND_LFI    32'h000002c8
`define DCMAC__C33_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C33_CTL_TX_SEND_RFI    32'h000002c9
`define DCMAC__C33_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C34_CTL_RX_CHECK_PREAMBLE    32'h000002ca
`define DCMAC__C34_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C34_CTL_RX_CHECK_SFD    32'h000002cb
`define DCMAC__C34_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C34_CTL_RX_DELETE_FCS    32'h000002cc
`define DCMAC__C34_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C34_CTL_RX_IGNORE_FCS    32'h000002cd
`define DCMAC__C34_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C34_CTL_RX_IGNORE_INRANGE    32'h000002ce
`define DCMAC__C34_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C34_CTL_RX_IS_CLAUSE_49    32'h000002cf
`define DCMAC__C34_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C34_CTL_RX_MAX_PACKET_LEN    32'h000002d0
`define DCMAC__C34_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C34_CTL_RX_PROCESS_LFI    32'h000002d1
`define DCMAC__C34_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C34_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002d2
`define DCMAC__C34_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C34_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002d3
`define DCMAC__C34_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C34_CTL_TX_FCS_INS_ENABLE    32'h000002d4
`define DCMAC__C34_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C34_CTL_TX_IGNORE_FCS    32'h000002d5
`define DCMAC__C34_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C34_CTL_TX_IPG_VALUE    32'h000002d6
`define DCMAC__C34_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C34_CTL_TX_SEND_IDLE    32'h000002d7
`define DCMAC__C34_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C34_CTL_TX_SEND_LFI    32'h000002d8
`define DCMAC__C34_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C34_CTL_TX_SEND_RFI    32'h000002d9
`define DCMAC__C34_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C35_CTL_RX_CHECK_PREAMBLE    32'h000002da
`define DCMAC__C35_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C35_CTL_RX_CHECK_SFD    32'h000002db
`define DCMAC__C35_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C35_CTL_RX_DELETE_FCS    32'h000002dc
`define DCMAC__C35_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C35_CTL_RX_IGNORE_FCS    32'h000002dd
`define DCMAC__C35_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C35_CTL_RX_IGNORE_INRANGE    32'h000002de
`define DCMAC__C35_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C35_CTL_RX_IS_CLAUSE_49    32'h000002df
`define DCMAC__C35_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C35_CTL_RX_MAX_PACKET_LEN    32'h000002e0
`define DCMAC__C35_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C35_CTL_RX_PROCESS_LFI    32'h000002e1
`define DCMAC__C35_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C35_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002e2
`define DCMAC__C35_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C35_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002e3
`define DCMAC__C35_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C35_CTL_TX_FCS_INS_ENABLE    32'h000002e4
`define DCMAC__C35_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C35_CTL_TX_IGNORE_FCS    32'h000002e5
`define DCMAC__C35_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C35_CTL_TX_IPG_VALUE    32'h000002e6
`define DCMAC__C35_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C35_CTL_TX_SEND_IDLE    32'h000002e7
`define DCMAC__C35_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C35_CTL_TX_SEND_LFI    32'h000002e8
`define DCMAC__C35_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C35_CTL_TX_SEND_RFI    32'h000002e9
`define DCMAC__C35_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C36_CTL_RX_CHECK_PREAMBLE    32'h000002ea
`define DCMAC__C36_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C36_CTL_RX_CHECK_SFD    32'h000002eb
`define DCMAC__C36_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C36_CTL_RX_DELETE_FCS    32'h000002ec
`define DCMAC__C36_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C36_CTL_RX_IGNORE_FCS    32'h000002ed
`define DCMAC__C36_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C36_CTL_RX_IGNORE_INRANGE    32'h000002ee
`define DCMAC__C36_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C36_CTL_RX_IS_CLAUSE_49    32'h000002ef
`define DCMAC__C36_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C36_CTL_RX_MAX_PACKET_LEN    32'h000002f0
`define DCMAC__C36_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C36_CTL_RX_PROCESS_LFI    32'h000002f1
`define DCMAC__C36_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C36_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000002f2
`define DCMAC__C36_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C36_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000002f3
`define DCMAC__C36_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C36_CTL_TX_FCS_INS_ENABLE    32'h000002f4
`define DCMAC__C36_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C36_CTL_TX_IGNORE_FCS    32'h000002f5
`define DCMAC__C36_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C36_CTL_TX_IPG_VALUE    32'h000002f6
`define DCMAC__C36_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C36_CTL_TX_SEND_IDLE    32'h000002f7
`define DCMAC__C36_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C36_CTL_TX_SEND_LFI    32'h000002f8
`define DCMAC__C36_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C36_CTL_TX_SEND_RFI    32'h000002f9
`define DCMAC__C36_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C37_CTL_RX_CHECK_PREAMBLE    32'h000002fa
`define DCMAC__C37_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C37_CTL_RX_CHECK_SFD    32'h000002fb
`define DCMAC__C37_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C37_CTL_RX_DELETE_FCS    32'h000002fc
`define DCMAC__C37_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C37_CTL_RX_IGNORE_FCS    32'h000002fd
`define DCMAC__C37_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C37_CTL_RX_IGNORE_INRANGE    32'h000002fe
`define DCMAC__C37_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C37_CTL_RX_IS_CLAUSE_49    32'h000002ff
`define DCMAC__C37_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C37_CTL_RX_MAX_PACKET_LEN    32'h00000300
`define DCMAC__C37_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C37_CTL_RX_PROCESS_LFI    32'h00000301
`define DCMAC__C37_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C37_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000302
`define DCMAC__C37_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C37_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000303
`define DCMAC__C37_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C37_CTL_TX_FCS_INS_ENABLE    32'h00000304
`define DCMAC__C37_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C37_CTL_TX_IGNORE_FCS    32'h00000305
`define DCMAC__C37_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C37_CTL_TX_IPG_VALUE    32'h00000306
`define DCMAC__C37_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C37_CTL_TX_SEND_IDLE    32'h00000307
`define DCMAC__C37_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C37_CTL_TX_SEND_LFI    32'h00000308
`define DCMAC__C37_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C37_CTL_TX_SEND_RFI    32'h00000309
`define DCMAC__C37_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C38_CTL_RX_CHECK_PREAMBLE    32'h0000030a
`define DCMAC__C38_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C38_CTL_RX_CHECK_SFD    32'h0000030b
`define DCMAC__C38_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C38_CTL_RX_DELETE_FCS    32'h0000030c
`define DCMAC__C38_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C38_CTL_RX_IGNORE_FCS    32'h0000030d
`define DCMAC__C38_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C38_CTL_RX_IGNORE_INRANGE    32'h0000030e
`define DCMAC__C38_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C38_CTL_RX_IS_CLAUSE_49    32'h0000030f
`define DCMAC__C38_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C38_CTL_RX_MAX_PACKET_LEN    32'h00000310
`define DCMAC__C38_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C38_CTL_RX_PROCESS_LFI    32'h00000311
`define DCMAC__C38_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C38_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000312
`define DCMAC__C38_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C38_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000313
`define DCMAC__C38_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C38_CTL_TX_FCS_INS_ENABLE    32'h00000314
`define DCMAC__C38_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C38_CTL_TX_IGNORE_FCS    32'h00000315
`define DCMAC__C38_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C38_CTL_TX_IPG_VALUE    32'h00000316
`define DCMAC__C38_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C38_CTL_TX_SEND_IDLE    32'h00000317
`define DCMAC__C38_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C38_CTL_TX_SEND_LFI    32'h00000318
`define DCMAC__C38_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C38_CTL_TX_SEND_RFI    32'h00000319
`define DCMAC__C38_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C39_CTL_RX_CHECK_PREAMBLE    32'h0000031a
`define DCMAC__C39_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C39_CTL_RX_CHECK_SFD    32'h0000031b
`define DCMAC__C39_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C39_CTL_RX_DELETE_FCS    32'h0000031c
`define DCMAC__C39_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C39_CTL_RX_IGNORE_FCS    32'h0000031d
`define DCMAC__C39_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C39_CTL_RX_IGNORE_INRANGE    32'h0000031e
`define DCMAC__C39_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C39_CTL_RX_IS_CLAUSE_49    32'h0000031f
`define DCMAC__C39_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C39_CTL_RX_MAX_PACKET_LEN    32'h00000320
`define DCMAC__C39_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C39_CTL_RX_PROCESS_LFI    32'h00000321
`define DCMAC__C39_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C39_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000322
`define DCMAC__C39_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C39_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000323
`define DCMAC__C39_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C39_CTL_TX_FCS_INS_ENABLE    32'h00000324
`define DCMAC__C39_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C39_CTL_TX_IGNORE_FCS    32'h00000325
`define DCMAC__C39_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C39_CTL_TX_IPG_VALUE    32'h00000326
`define DCMAC__C39_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C39_CTL_TX_SEND_IDLE    32'h00000327
`define DCMAC__C39_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C39_CTL_TX_SEND_LFI    32'h00000328
`define DCMAC__C39_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C39_CTL_TX_SEND_RFI    32'h00000329
`define DCMAC__C39_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C3_CTL_PCS_RX_TS_EN    32'h0000032a
`define DCMAC__C3_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_ACK    32'h0000032b
`define DCMAC__C3_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_ETYPE_GCP    32'h0000032c
`define DCMAC__C3_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_ETYPE_GPP    32'h0000032d
`define DCMAC__C3_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_ETYPE_PCP    32'h0000032e
`define DCMAC__C3_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_ETYPE_PPP    32'h0000032f
`define DCMAC__C3_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_MCAST_GCP    32'h00000330
`define DCMAC__C3_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_MCAST_GPP    32'h00000331
`define DCMAC__C3_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_MCAST_PCP    32'h00000332
`define DCMAC__C3_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_MCAST_PPP    32'h00000333
`define DCMAC__C3_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_OPCODE_GCP    32'h00000334
`define DCMAC__C3_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_OPCODE_GPP    32'h00000335
`define DCMAC__C3_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_OPCODE_PCP    32'h00000336
`define DCMAC__C3_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_OPCODE_PPP    32'h00000337
`define DCMAC__C3_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_PREAMBLE    32'h00000338
`define DCMAC__C3_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_SA_GCP    32'h00000339
`define DCMAC__C3_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_SA_GPP    32'h0000033a
`define DCMAC__C3_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_SA_PCP    32'h0000033b
`define DCMAC__C3_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_SA_PPP    32'h0000033c
`define DCMAC__C3_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_SFD    32'h0000033d
`define DCMAC__C3_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_UCAST_GCP    32'h0000033e
`define DCMAC__C3_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_UCAST_GPP    32'h0000033f
`define DCMAC__C3_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_UCAST_PCP    32'h00000340
`define DCMAC__C3_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C3_CTL_RX_CHECK_UCAST_PPP    32'h00000341
`define DCMAC__C3_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C3_CTL_RX_DEGRADE_ACT_THRESH    32'h00000342
`define DCMAC__C3_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C3_CTL_RX_DEGRADE_DEACT_THRESH    32'h00000343
`define DCMAC__C3_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C3_CTL_RX_DEGRADE_ENABLE    32'h00000344
`define DCMAC__C3_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C3_CTL_RX_DEGRADE_INTERVAL    32'h00000345
`define DCMAC__C3_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C3_CTL_RX_DELETE_FCS    32'h00000346
`define DCMAC__C3_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C3_CTL_RX_ENABLE_GCP    32'h00000347
`define DCMAC__C3_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C3_CTL_RX_ENABLE_GPP    32'h00000348
`define DCMAC__C3_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C3_CTL_RX_ENABLE_PCP    32'h00000349
`define DCMAC__C3_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C3_CTL_RX_ENABLE_PPP    32'h0000034a
`define DCMAC__C3_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C3_CTL_RX_ETYPE_GCP    32'h0000034b
`define DCMAC__C3_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C3_CTL_RX_ETYPE_GPP    32'h0000034c
`define DCMAC__C3_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C3_CTL_RX_ETYPE_PCP    32'h0000034d
`define DCMAC__C3_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C3_CTL_RX_ETYPE_PPP    32'h0000034e
`define DCMAC__C3_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C3_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h0000034f
`define DCMAC__C3_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C3_CTL_RX_FEC_BYPASS_CORRECTION    32'h00000350
`define DCMAC__C3_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C3_CTL_RX_FEC_BYPASS_INDICATION    32'h00000351
`define DCMAC__C3_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C3_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h00000352
`define DCMAC__C3_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C3_CTL_RX_FEC_MODE    32'h00000353
`define DCMAC__C3_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C3_CTL_RX_FEC_TRANSCODE_BYPASS    32'h00000354
`define DCMAC__C3_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C3_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h00000355
`define DCMAC__C3_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C3_CTL_RX_FLEXIF_PCS_WIDE_MODE    32'h00000356
`define DCMAC__C3_CTL_RX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C3_CTL_RX_FLEXIF_SELECT    32'h00000357
`define DCMAC__C3_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C3_CTL_RX_FORWARD_CONTROL    32'h00000358
`define DCMAC__C3_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C3_CTL_RX_IGNORE_FCS    32'h00000359
`define DCMAC__C3_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C3_CTL_RX_IGNORE_INRANGE    32'h0000035a
`define DCMAC__C3_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C3_CTL_RX_IS_CLAUSE_49    32'h0000035b
`define DCMAC__C3_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C3_CTL_RX_MAX_PACKET_LEN    32'h0000035c
`define DCMAC__C3_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C3_CTL_RX_OPCODE_GPP    32'h0000035d
`define DCMAC__C3_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C3_CTL_RX_OPCODE_MAX_GCP    32'h0000035e
`define DCMAC__C3_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C3_CTL_RX_OPCODE_MAX_PCP    32'h0000035f
`define DCMAC__C3_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C3_CTL_RX_OPCODE_MIN_GCP    32'h00000360
`define DCMAC__C3_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C3_CTL_RX_OPCODE_MIN_PCP    32'h00000361
`define DCMAC__C3_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C3_CTL_RX_OPCODE_PPP    32'h00000362
`define DCMAC__C3_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C3_CTL_RX_PAUSE_DA_MCAST    32'h00000363
`define DCMAC__C3_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C3_CTL_RX_PAUSE_DA_UCAST    32'h00000364
`define DCMAC__C3_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C3_CTL_RX_PAUSE_SA    32'h00000365
`define DCMAC__C3_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C3_CTL_RX_PMA_LANE_MUX    32'h00000366
`define DCMAC__C3_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C3_CTL_RX_PROCESS_LFI    32'h00000367
`define DCMAC__C3_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C3_CTL_RX_PTP_LATENCY_ADJUST    32'h00000368
`define DCMAC__C3_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C3_CTL_RX_PTP_ST_OFFSET    32'h00000369
`define DCMAC__C3_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C3_CTL_RX_TEST_PATTERN    32'h0000036a
`define DCMAC__C3_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C3_CTL_RX_TICK_REG_MODE_SEL    32'h0000036b
`define DCMAC__C3_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C3_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h0000036c
`define DCMAC__C3_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C3_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h0000036d
`define DCMAC__C3_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C3_CTL_TX_CORRUPT_FCS_ON_ERR    32'h0000036e
`define DCMAC__C3_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C3_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h0000036f
`define DCMAC__C3_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C3_CTL_TX_DA_GPP    32'h00000370
`define DCMAC__C3_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C3_CTL_TX_DA_PPP    32'h00000371
`define DCMAC__C3_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C3_CTL_TX_ETHERTYPE_GPP    32'h00000372
`define DCMAC__C3_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C3_CTL_TX_ETHERTYPE_PPP    32'h00000373
`define DCMAC__C3_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C3_CTL_TX_FCS_INS_ENABLE    32'h00000374
`define DCMAC__C3_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C3_CTL_TX_FEC_FOUR_LANE_PMD    32'h00000375
`define DCMAC__C3_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C3_CTL_TX_FEC_MODE    32'h00000376
`define DCMAC__C3_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C3_CTL_TX_FEC_TRANSCODE_BYPASS    32'h00000377
`define DCMAC__C3_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C3_CTL_TX_FLEXIF_AM_MODE    32'h00000378
`define DCMAC__C3_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C3_CTL_TX_FLEXIF_PCS_WIDE_MODE    32'h00000379
`define DCMAC__C3_CTL_TX_FLEXIF_PCS_WIDE_MODE_SZ 40

`define DCMAC__C3_CTL_TX_FLEXIF_SELECT    32'h0000037a
`define DCMAC__C3_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C3_CTL_TX_IGNORE_FCS    32'h0000037b
`define DCMAC__C3_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C3_CTL_TX_IPG_VALUE    32'h0000037c
`define DCMAC__C3_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C3_CTL_TX_OPCODE_GPP    32'h0000037d
`define DCMAC__C3_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C3_CTL_TX_OPCODE_PPP    32'h0000037e
`define DCMAC__C3_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA0    32'h0000037f
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA1    32'h00000380
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA2    32'h00000381
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA3    32'h00000382
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA4    32'h00000383
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA5    32'h00000384
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA6    32'h00000385
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA7    32'h00000386
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_QUANTA8    32'h00000387
`define DCMAC__C3_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C3_CTL_TX_PAUSE_REFRESH_TIMER    32'h00000388
`define DCMAC__C3_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C3_CTL_TX_PMA_LANE_MUX    32'h00000389
`define DCMAC__C3_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C3_CTL_TX_PTP_1STEP_ENABLE    32'h0000038a
`define DCMAC__C3_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C3_CTL_TX_PTP_LATENCY_ADJUST    32'h0000038b
`define DCMAC__C3_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C3_CTL_TX_PTP_SAT_ENABLE    32'h0000038c
`define DCMAC__C3_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C3_CTL_TX_PTP_ST_OFFSET    32'h0000038d
`define DCMAC__C3_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C3_CTL_TX_SA_GPP    32'h0000038e
`define DCMAC__C3_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C3_CTL_TX_SA_PPP    32'h0000038f
`define DCMAC__C3_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C3_CTL_TX_SEND_IDLE    32'h00000390
`define DCMAC__C3_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C3_CTL_TX_SEND_LFI    32'h00000391
`define DCMAC__C3_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C3_CTL_TX_SEND_RFI    32'h00000392
`define DCMAC__C3_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C3_CTL_TX_TICK_REG_MODE_SEL    32'h00000393
`define DCMAC__C3_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C3_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000394
`define DCMAC__C3_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C3_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h00000395
`define DCMAC__C3_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C4_CTL_PCS_RX_TS_EN    32'h00000396
`define DCMAC__C4_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_ACK    32'h00000397
`define DCMAC__C4_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_ETYPE_GCP    32'h00000398
`define DCMAC__C4_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_ETYPE_GPP    32'h00000399
`define DCMAC__C4_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_ETYPE_PCP    32'h0000039a
`define DCMAC__C4_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_ETYPE_PPP    32'h0000039b
`define DCMAC__C4_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_MCAST_GCP    32'h0000039c
`define DCMAC__C4_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_MCAST_GPP    32'h0000039d
`define DCMAC__C4_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_MCAST_PCP    32'h0000039e
`define DCMAC__C4_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_MCAST_PPP    32'h0000039f
`define DCMAC__C4_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_OPCODE_GCP    32'h000003a0
`define DCMAC__C4_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_OPCODE_GPP    32'h000003a1
`define DCMAC__C4_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_OPCODE_PCP    32'h000003a2
`define DCMAC__C4_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_OPCODE_PPP    32'h000003a3
`define DCMAC__C4_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_PREAMBLE    32'h000003a4
`define DCMAC__C4_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_SA_GCP    32'h000003a5
`define DCMAC__C4_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_SA_GPP    32'h000003a6
`define DCMAC__C4_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_SA_PCP    32'h000003a7
`define DCMAC__C4_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_SA_PPP    32'h000003a8
`define DCMAC__C4_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_SFD    32'h000003a9
`define DCMAC__C4_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_UCAST_GCP    32'h000003aa
`define DCMAC__C4_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_UCAST_GPP    32'h000003ab
`define DCMAC__C4_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_UCAST_PCP    32'h000003ac
`define DCMAC__C4_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C4_CTL_RX_CHECK_UCAST_PPP    32'h000003ad
`define DCMAC__C4_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C4_CTL_RX_DATA_RATE    32'h000003ae
`define DCMAC__C4_CTL_RX_DATA_RATE_SZ 1

`define DCMAC__C4_CTL_RX_DEGRADE_ACT_THRESH    32'h000003af
`define DCMAC__C4_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C4_CTL_RX_DEGRADE_DEACT_THRESH    32'h000003b0
`define DCMAC__C4_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C4_CTL_RX_DEGRADE_ENABLE    32'h000003b1
`define DCMAC__C4_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C4_CTL_RX_DEGRADE_INTERVAL    32'h000003b2
`define DCMAC__C4_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C4_CTL_RX_DELETE_FCS    32'h000003b3
`define DCMAC__C4_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C4_CTL_RX_ENABLE_GCP    32'h000003b4
`define DCMAC__C4_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C4_CTL_RX_ENABLE_GPP    32'h000003b5
`define DCMAC__C4_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C4_CTL_RX_ENABLE_PCP    32'h000003b6
`define DCMAC__C4_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C4_CTL_RX_ENABLE_PPP    32'h000003b7
`define DCMAC__C4_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C4_CTL_RX_ETYPE_GCP    32'h000003b8
`define DCMAC__C4_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C4_CTL_RX_ETYPE_GPP    32'h000003b9
`define DCMAC__C4_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C4_CTL_RX_ETYPE_PCP    32'h000003ba
`define DCMAC__C4_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C4_CTL_RX_ETYPE_PPP    32'h000003bb
`define DCMAC__C4_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C4_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h000003bc
`define DCMAC__C4_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C4_CTL_RX_FEC_BYPASS_CORRECTION    32'h000003bd
`define DCMAC__C4_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C4_CTL_RX_FEC_BYPASS_INDICATION    32'h000003be
`define DCMAC__C4_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C4_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h000003bf
`define DCMAC__C4_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C4_CTL_RX_FEC_MODE    32'h000003c0
`define DCMAC__C4_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C4_CTL_RX_FEC_TRANSCODE_BYPASS    32'h000003c1
`define DCMAC__C4_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C4_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h000003c2
`define DCMAC__C4_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C4_CTL_RX_FLEXIF_SELECT    32'h000003c3
`define DCMAC__C4_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C4_CTL_RX_FORWARD_CONTROL    32'h000003c4
`define DCMAC__C4_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C4_CTL_RX_IGNORE_FCS    32'h000003c5
`define DCMAC__C4_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C4_CTL_RX_IGNORE_INRANGE    32'h000003c6
`define DCMAC__C4_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C4_CTL_RX_IS_CLAUSE_49    32'h000003c7
`define DCMAC__C4_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C4_CTL_RX_MAX_PACKET_LEN    32'h000003c8
`define DCMAC__C4_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C4_CTL_RX_OPCODE_GPP    32'h000003c9
`define DCMAC__C4_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C4_CTL_RX_OPCODE_MAX_GCP    32'h000003ca
`define DCMAC__C4_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C4_CTL_RX_OPCODE_MAX_PCP    32'h000003cb
`define DCMAC__C4_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C4_CTL_RX_OPCODE_MIN_GCP    32'h000003cc
`define DCMAC__C4_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C4_CTL_RX_OPCODE_MIN_PCP    32'h000003cd
`define DCMAC__C4_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C4_CTL_RX_OPCODE_PPP    32'h000003ce
`define DCMAC__C4_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C4_CTL_RX_PAUSE_DA_MCAST    32'h000003cf
`define DCMAC__C4_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C4_CTL_RX_PAUSE_DA_UCAST    32'h000003d0
`define DCMAC__C4_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C4_CTL_RX_PAUSE_SA    32'h000003d1
`define DCMAC__C4_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C4_CTL_RX_PMA_LANE_MUX    32'h000003d2
`define DCMAC__C4_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C4_CTL_RX_PROCESS_LFI    32'h000003d3
`define DCMAC__C4_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C4_CTL_RX_PTP_LATENCY_ADJUST    32'h000003d4
`define DCMAC__C4_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C4_CTL_RX_PTP_ST_OFFSET    32'h000003d5
`define DCMAC__C4_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C4_CTL_RX_TEST_PATTERN    32'h000003d6
`define DCMAC__C4_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C4_CTL_RX_TICK_REG_MODE_SEL    32'h000003d7
`define DCMAC__C4_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C4_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h000003d8
`define DCMAC__C4_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C4_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h000003d9
`define DCMAC__C4_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C4_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE    32'h000003da
`define DCMAC__C4_CTL_TX_ALT_SERDES_CLK_MUX_DISABLE_SZ 40

`define DCMAC__C4_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000003db
`define DCMAC__C4_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C4_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000003dc
`define DCMAC__C4_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C4_CTL_TX_DATA_RATE    32'h000003dd
`define DCMAC__C4_CTL_TX_DATA_RATE_SZ 1

`define DCMAC__C4_CTL_TX_DA_GPP    32'h000003de
`define DCMAC__C4_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C4_CTL_TX_DA_PPP    32'h000003df
`define DCMAC__C4_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C4_CTL_TX_ETHERTYPE_GPP    32'h000003e0
`define DCMAC__C4_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C4_CTL_TX_ETHERTYPE_PPP    32'h000003e1
`define DCMAC__C4_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C4_CTL_TX_FCS_INS_ENABLE    32'h000003e2
`define DCMAC__C4_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C4_CTL_TX_FEC_FOUR_LANE_PMD    32'h000003e3
`define DCMAC__C4_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C4_CTL_TX_FEC_MODE    32'h000003e4
`define DCMAC__C4_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C4_CTL_TX_FEC_TRANSCODE_BYPASS    32'h000003e5
`define DCMAC__C4_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C4_CTL_TX_FLEXIF_AM_MODE    32'h000003e6
`define DCMAC__C4_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C4_CTL_TX_FLEXIF_SELECT    32'h000003e7
`define DCMAC__C4_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C4_CTL_TX_IGNORE_FCS    32'h000003e8
`define DCMAC__C4_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C4_CTL_TX_IPG_VALUE    32'h000003e9
`define DCMAC__C4_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C4_CTL_TX_OPCODE_GPP    32'h000003ea
`define DCMAC__C4_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C4_CTL_TX_OPCODE_PPP    32'h000003eb
`define DCMAC__C4_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA0    32'h000003ec
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA1    32'h000003ed
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA2    32'h000003ee
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA3    32'h000003ef
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA4    32'h000003f0
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA5    32'h000003f1
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA6    32'h000003f2
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA7    32'h000003f3
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_QUANTA8    32'h000003f4
`define DCMAC__C4_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C4_CTL_TX_PAUSE_REFRESH_TIMER    32'h000003f5
`define DCMAC__C4_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C4_CTL_TX_PMA_LANE_MUX    32'h000003f6
`define DCMAC__C4_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C4_CTL_TX_PTP_1STEP_ENABLE    32'h000003f7
`define DCMAC__C4_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C4_CTL_TX_PTP_LATENCY_ADJUST    32'h000003f8
`define DCMAC__C4_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C4_CTL_TX_PTP_SAT_ENABLE    32'h000003f9
`define DCMAC__C4_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C4_CTL_TX_PTP_ST_OFFSET    32'h000003fa
`define DCMAC__C4_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C4_CTL_TX_SA_GPP    32'h000003fb
`define DCMAC__C4_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C4_CTL_TX_SA_PPP    32'h000003fc
`define DCMAC__C4_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C4_CTL_TX_SEND_IDLE    32'h000003fd
`define DCMAC__C4_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C4_CTL_TX_SEND_LFI    32'h000003fe
`define DCMAC__C4_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C4_CTL_TX_SEND_RFI    32'h000003ff
`define DCMAC__C4_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C4_CTL_TX_TICK_REG_MODE_SEL    32'h00000400
`define DCMAC__C4_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C4_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000401
`define DCMAC__C4_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C4_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h00000402
`define DCMAC__C4_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C5_CTL_PCS_RX_TS_EN    32'h00000403
`define DCMAC__C5_CTL_PCS_RX_TS_EN_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_ACK    32'h00000404
`define DCMAC__C5_CTL_RX_CHECK_ACK_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_ETYPE_GCP    32'h00000405
`define DCMAC__C5_CTL_RX_CHECK_ETYPE_GCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_ETYPE_GPP    32'h00000406
`define DCMAC__C5_CTL_RX_CHECK_ETYPE_GPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_ETYPE_PCP    32'h00000407
`define DCMAC__C5_CTL_RX_CHECK_ETYPE_PCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_ETYPE_PPP    32'h00000408
`define DCMAC__C5_CTL_RX_CHECK_ETYPE_PPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_MCAST_GCP    32'h00000409
`define DCMAC__C5_CTL_RX_CHECK_MCAST_GCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_MCAST_GPP    32'h0000040a
`define DCMAC__C5_CTL_RX_CHECK_MCAST_GPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_MCAST_PCP    32'h0000040b
`define DCMAC__C5_CTL_RX_CHECK_MCAST_PCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_MCAST_PPP    32'h0000040c
`define DCMAC__C5_CTL_RX_CHECK_MCAST_PPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_OPCODE_GCP    32'h0000040d
`define DCMAC__C5_CTL_RX_CHECK_OPCODE_GCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_OPCODE_GPP    32'h0000040e
`define DCMAC__C5_CTL_RX_CHECK_OPCODE_GPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_OPCODE_PCP    32'h0000040f
`define DCMAC__C5_CTL_RX_CHECK_OPCODE_PCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_OPCODE_PPP    32'h00000410
`define DCMAC__C5_CTL_RX_CHECK_OPCODE_PPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_PREAMBLE    32'h00000411
`define DCMAC__C5_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_SA_GCP    32'h00000412
`define DCMAC__C5_CTL_RX_CHECK_SA_GCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_SA_GPP    32'h00000413
`define DCMAC__C5_CTL_RX_CHECK_SA_GPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_SA_PCP    32'h00000414
`define DCMAC__C5_CTL_RX_CHECK_SA_PCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_SA_PPP    32'h00000415
`define DCMAC__C5_CTL_RX_CHECK_SA_PPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_SFD    32'h00000416
`define DCMAC__C5_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_UCAST_GCP    32'h00000417
`define DCMAC__C5_CTL_RX_CHECK_UCAST_GCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_UCAST_GPP    32'h00000418
`define DCMAC__C5_CTL_RX_CHECK_UCAST_GPP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_UCAST_PCP    32'h00000419
`define DCMAC__C5_CTL_RX_CHECK_UCAST_PCP_SZ 40

`define DCMAC__C5_CTL_RX_CHECK_UCAST_PPP    32'h0000041a
`define DCMAC__C5_CTL_RX_CHECK_UCAST_PPP_SZ 40

`define DCMAC__C5_CTL_RX_DEGRADE_ACT_THRESH    32'h0000041b
`define DCMAC__C5_CTL_RX_DEGRADE_ACT_THRESH_SZ 32

`define DCMAC__C5_CTL_RX_DEGRADE_DEACT_THRESH    32'h0000041c
`define DCMAC__C5_CTL_RX_DEGRADE_DEACT_THRESH_SZ 32

`define DCMAC__C5_CTL_RX_DEGRADE_ENABLE    32'h0000041d
`define DCMAC__C5_CTL_RX_DEGRADE_ENABLE_SZ 40

`define DCMAC__C5_CTL_RX_DEGRADE_INTERVAL    32'h0000041e
`define DCMAC__C5_CTL_RX_DEGRADE_INTERVAL_SZ 32

`define DCMAC__C5_CTL_RX_DELETE_FCS    32'h0000041f
`define DCMAC__C5_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C5_CTL_RX_ENABLE_GCP    32'h00000420
`define DCMAC__C5_CTL_RX_ENABLE_GCP_SZ 40

`define DCMAC__C5_CTL_RX_ENABLE_GPP    32'h00000421
`define DCMAC__C5_CTL_RX_ENABLE_GPP_SZ 40

`define DCMAC__C5_CTL_RX_ENABLE_PCP    32'h00000422
`define DCMAC__C5_CTL_RX_ENABLE_PCP_SZ 40

`define DCMAC__C5_CTL_RX_ENABLE_PPP    32'h00000423
`define DCMAC__C5_CTL_RX_ENABLE_PPP_SZ 40

`define DCMAC__C5_CTL_RX_ETYPE_GCP    32'h00000424
`define DCMAC__C5_CTL_RX_ETYPE_GCP_SZ 16

`define DCMAC__C5_CTL_RX_ETYPE_GPP    32'h00000425
`define DCMAC__C5_CTL_RX_ETYPE_GPP_SZ 16

`define DCMAC__C5_CTL_RX_ETYPE_PCP    32'h00000426
`define DCMAC__C5_CTL_RX_ETYPE_PCP_SZ 16

`define DCMAC__C5_CTL_RX_ETYPE_PPP    32'h00000427
`define DCMAC__C5_CTL_RX_ETYPE_PPP_SZ 16

`define DCMAC__C5_CTL_RX_FEC_ALIGNMENT_BYPASS    32'h00000428
`define DCMAC__C5_CTL_RX_FEC_ALIGNMENT_BYPASS_SZ 40

`define DCMAC__C5_CTL_RX_FEC_BYPASS_CORRECTION    32'h00000429
`define DCMAC__C5_CTL_RX_FEC_BYPASS_CORRECTION_SZ 40

`define DCMAC__C5_CTL_RX_FEC_BYPASS_INDICATION    32'h0000042a
`define DCMAC__C5_CTL_RX_FEC_BYPASS_INDICATION_SZ 40

`define DCMAC__C5_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE    32'h0000042b
`define DCMAC__C5_CTL_RX_FEC_EXT_ALIGN_BUFF_ENABLE_SZ 40

`define DCMAC__C5_CTL_RX_FEC_MODE    32'h0000042c
`define DCMAC__C5_CTL_RX_FEC_MODE_SZ 5

`define DCMAC__C5_CTL_RX_FEC_TRANSCODE_BYPASS    32'h0000042d
`define DCMAC__C5_CTL_RX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C5_CTL_RX_FEC_TRANSCODE_CLAUSE49    32'h0000042e
`define DCMAC__C5_CTL_RX_FEC_TRANSCODE_CLAUSE49_SZ 40

`define DCMAC__C5_CTL_RX_FLEXIF_SELECT    32'h0000042f
`define DCMAC__C5_CTL_RX_FLEXIF_SELECT_SZ 2

`define DCMAC__C5_CTL_RX_FORWARD_CONTROL    32'h00000430
`define DCMAC__C5_CTL_RX_FORWARD_CONTROL_SZ 40

`define DCMAC__C5_CTL_RX_IGNORE_FCS    32'h00000431
`define DCMAC__C5_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C5_CTL_RX_IGNORE_INRANGE    32'h00000432
`define DCMAC__C5_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C5_CTL_RX_IS_CLAUSE_49    32'h00000433
`define DCMAC__C5_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C5_CTL_RX_MAX_PACKET_LEN    32'h00000434
`define DCMAC__C5_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C5_CTL_RX_OPCODE_GPP    32'h00000435
`define DCMAC__C5_CTL_RX_OPCODE_GPP_SZ 16

`define DCMAC__C5_CTL_RX_OPCODE_MAX_GCP    32'h00000436
`define DCMAC__C5_CTL_RX_OPCODE_MAX_GCP_SZ 16

`define DCMAC__C5_CTL_RX_OPCODE_MAX_PCP    32'h00000437
`define DCMAC__C5_CTL_RX_OPCODE_MAX_PCP_SZ 16

`define DCMAC__C5_CTL_RX_OPCODE_MIN_GCP    32'h00000438
`define DCMAC__C5_CTL_RX_OPCODE_MIN_GCP_SZ 16

`define DCMAC__C5_CTL_RX_OPCODE_MIN_PCP    32'h00000439
`define DCMAC__C5_CTL_RX_OPCODE_MIN_PCP_SZ 16

`define DCMAC__C5_CTL_RX_OPCODE_PPP    32'h0000043a
`define DCMAC__C5_CTL_RX_OPCODE_PPP_SZ 16

`define DCMAC__C5_CTL_RX_PAUSE_DA_MCAST    32'h0000043b
`define DCMAC__C5_CTL_RX_PAUSE_DA_MCAST_SZ 48

`define DCMAC__C5_CTL_RX_PAUSE_DA_UCAST    32'h0000043c
`define DCMAC__C5_CTL_RX_PAUSE_DA_UCAST_SZ 48

`define DCMAC__C5_CTL_RX_PAUSE_SA    32'h0000043d
`define DCMAC__C5_CTL_RX_PAUSE_SA_SZ 48

`define DCMAC__C5_CTL_RX_PMA_LANE_MUX    32'h0000043e
`define DCMAC__C5_CTL_RX_PMA_LANE_MUX_SZ 2

`define DCMAC__C5_CTL_RX_PROCESS_LFI    32'h0000043f
`define DCMAC__C5_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C5_CTL_RX_PTP_LATENCY_ADJUST    32'h00000440
`define DCMAC__C5_CTL_RX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C5_CTL_RX_PTP_ST_OFFSET    32'h00000441
`define DCMAC__C5_CTL_RX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C5_CTL_RX_TEST_PATTERN    32'h00000442
`define DCMAC__C5_CTL_RX_TEST_PATTERN_SZ 40

`define DCMAC__C5_CTL_RX_TICK_REG_MODE_SEL    32'h00000443
`define DCMAC__C5_CTL_RX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C5_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h00000444
`define DCMAC__C5_CTL_RX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C5_CTL_RX_USE_CUSTOM_VL_MARKER_IDS    32'h00000445
`define DCMAC__C5_CTL_RX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C5_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000446
`define DCMAC__C5_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C5_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000447
`define DCMAC__C5_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C5_CTL_TX_DA_GPP    32'h00000448
`define DCMAC__C5_CTL_TX_DA_GPP_SZ 48

`define DCMAC__C5_CTL_TX_DA_PPP    32'h00000449
`define DCMAC__C5_CTL_TX_DA_PPP_SZ 48

`define DCMAC__C5_CTL_TX_ETHERTYPE_GPP    32'h0000044a
`define DCMAC__C5_CTL_TX_ETHERTYPE_GPP_SZ 16

`define DCMAC__C5_CTL_TX_ETHERTYPE_PPP    32'h0000044b
`define DCMAC__C5_CTL_TX_ETHERTYPE_PPP_SZ 16

`define DCMAC__C5_CTL_TX_FCS_INS_ENABLE    32'h0000044c
`define DCMAC__C5_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C5_CTL_TX_FEC_FOUR_LANE_PMD    32'h0000044d
`define DCMAC__C5_CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define DCMAC__C5_CTL_TX_FEC_MODE    32'h0000044e
`define DCMAC__C5_CTL_TX_FEC_MODE_SZ 5

`define DCMAC__C5_CTL_TX_FEC_TRANSCODE_BYPASS    32'h0000044f
`define DCMAC__C5_CTL_TX_FEC_TRANSCODE_BYPASS_SZ 40

`define DCMAC__C5_CTL_TX_FLEXIF_AM_MODE    32'h00000450
`define DCMAC__C5_CTL_TX_FLEXIF_AM_MODE_SZ 40

`define DCMAC__C5_CTL_TX_FLEXIF_SELECT    32'h00000451
`define DCMAC__C5_CTL_TX_FLEXIF_SELECT_SZ 2

`define DCMAC__C5_CTL_TX_IGNORE_FCS    32'h00000452
`define DCMAC__C5_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C5_CTL_TX_IPG_VALUE    32'h00000453
`define DCMAC__C5_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C5_CTL_TX_OPCODE_GPP    32'h00000454
`define DCMAC__C5_CTL_TX_OPCODE_GPP_SZ 16

`define DCMAC__C5_CTL_TX_OPCODE_PPP    32'h00000455
`define DCMAC__C5_CTL_TX_OPCODE_PPP_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA0    32'h00000456
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA0_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA1    32'h00000457
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA1_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA2    32'h00000458
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA2_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA3    32'h00000459
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA3_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA4    32'h0000045a
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA4_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA5    32'h0000045b
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA5_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA6    32'h0000045c
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA6_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA7    32'h0000045d
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA7_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_QUANTA8    32'h0000045e
`define DCMAC__C5_CTL_TX_PAUSE_QUANTA8_SZ 16

`define DCMAC__C5_CTL_TX_PAUSE_REFRESH_TIMER    32'h0000045f
`define DCMAC__C5_CTL_TX_PAUSE_REFRESH_TIMER_SZ 16

`define DCMAC__C5_CTL_TX_PMA_LANE_MUX    32'h00000460
`define DCMAC__C5_CTL_TX_PMA_LANE_MUX_SZ 2

`define DCMAC__C5_CTL_TX_PTP_1STEP_ENABLE    32'h00000461
`define DCMAC__C5_CTL_TX_PTP_1STEP_ENABLE_SZ 40

`define DCMAC__C5_CTL_TX_PTP_LATENCY_ADJUST    32'h00000462
`define DCMAC__C5_CTL_TX_PTP_LATENCY_ADJUST_SZ 20

`define DCMAC__C5_CTL_TX_PTP_SAT_ENABLE    32'h00000463
`define DCMAC__C5_CTL_TX_PTP_SAT_ENABLE_SZ 2

`define DCMAC__C5_CTL_TX_PTP_ST_OFFSET    32'h00000464
`define DCMAC__C5_CTL_TX_PTP_ST_OFFSET_SZ 16

`define DCMAC__C5_CTL_TX_SA_GPP    32'h00000465
`define DCMAC__C5_CTL_TX_SA_GPP_SZ 48

`define DCMAC__C5_CTL_TX_SA_PPP    32'h00000466
`define DCMAC__C5_CTL_TX_SA_PPP_SZ 48

`define DCMAC__C5_CTL_TX_SEND_IDLE    32'h00000467
`define DCMAC__C5_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C5_CTL_TX_SEND_LFI    32'h00000468
`define DCMAC__C5_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C5_CTL_TX_SEND_RFI    32'h00000469
`define DCMAC__C5_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C5_CTL_TX_TICK_REG_MODE_SEL    32'h0000046a
`define DCMAC__C5_CTL_TX_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__C5_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1    32'h0000046b
`define DCMAC__C5_CTL_TX_USE_CUSTOM_VL_LENGTH_MINUS1_SZ 40

`define DCMAC__C5_CTL_TX_USE_CUSTOM_VL_MARKER_IDS    32'h0000046c
`define DCMAC__C5_CTL_TX_USE_CUSTOM_VL_MARKER_IDS_SZ 40

`define DCMAC__C6_CTL_RX_CHECK_PREAMBLE    32'h0000046d
`define DCMAC__C6_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C6_CTL_RX_CHECK_SFD    32'h0000046e
`define DCMAC__C6_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C6_CTL_RX_DELETE_FCS    32'h0000046f
`define DCMAC__C6_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C6_CTL_RX_IGNORE_FCS    32'h00000470
`define DCMAC__C6_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C6_CTL_RX_IGNORE_INRANGE    32'h00000471
`define DCMAC__C6_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C6_CTL_RX_IS_CLAUSE_49    32'h00000472
`define DCMAC__C6_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C6_CTL_RX_MAX_PACKET_LEN    32'h00000473
`define DCMAC__C6_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C6_CTL_RX_PROCESS_LFI    32'h00000474
`define DCMAC__C6_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C6_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000475
`define DCMAC__C6_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C6_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000476
`define DCMAC__C6_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C6_CTL_TX_FCS_INS_ENABLE    32'h00000477
`define DCMAC__C6_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C6_CTL_TX_IGNORE_FCS    32'h00000478
`define DCMAC__C6_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C6_CTL_TX_IPG_VALUE    32'h00000479
`define DCMAC__C6_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C6_CTL_TX_SEND_IDLE    32'h0000047a
`define DCMAC__C6_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C6_CTL_TX_SEND_LFI    32'h0000047b
`define DCMAC__C6_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C6_CTL_TX_SEND_RFI    32'h0000047c
`define DCMAC__C6_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C7_CTL_RX_CHECK_PREAMBLE    32'h0000047d
`define DCMAC__C7_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C7_CTL_RX_CHECK_SFD    32'h0000047e
`define DCMAC__C7_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C7_CTL_RX_DELETE_FCS    32'h0000047f
`define DCMAC__C7_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C7_CTL_RX_IGNORE_FCS    32'h00000480
`define DCMAC__C7_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C7_CTL_RX_IGNORE_INRANGE    32'h00000481
`define DCMAC__C7_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C7_CTL_RX_IS_CLAUSE_49    32'h00000482
`define DCMAC__C7_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C7_CTL_RX_MAX_PACKET_LEN    32'h00000483
`define DCMAC__C7_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C7_CTL_RX_PROCESS_LFI    32'h00000484
`define DCMAC__C7_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C7_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000485
`define DCMAC__C7_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C7_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000486
`define DCMAC__C7_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C7_CTL_TX_FCS_INS_ENABLE    32'h00000487
`define DCMAC__C7_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C7_CTL_TX_IGNORE_FCS    32'h00000488
`define DCMAC__C7_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C7_CTL_TX_IPG_VALUE    32'h00000489
`define DCMAC__C7_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C7_CTL_TX_SEND_IDLE    32'h0000048a
`define DCMAC__C7_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C7_CTL_TX_SEND_LFI    32'h0000048b
`define DCMAC__C7_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C7_CTL_TX_SEND_RFI    32'h0000048c
`define DCMAC__C7_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C8_CTL_RX_CHECK_PREAMBLE    32'h0000048d
`define DCMAC__C8_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C8_CTL_RX_CHECK_SFD    32'h0000048e
`define DCMAC__C8_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C8_CTL_RX_DELETE_FCS    32'h0000048f
`define DCMAC__C8_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C8_CTL_RX_IGNORE_FCS    32'h00000490
`define DCMAC__C8_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C8_CTL_RX_IGNORE_INRANGE    32'h00000491
`define DCMAC__C8_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C8_CTL_RX_IS_CLAUSE_49    32'h00000492
`define DCMAC__C8_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C8_CTL_RX_MAX_PACKET_LEN    32'h00000493
`define DCMAC__C8_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C8_CTL_RX_PROCESS_LFI    32'h00000494
`define DCMAC__C8_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C8_CTL_TX_CORRUPT_FCS_ON_ERR    32'h00000495
`define DCMAC__C8_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C8_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h00000496
`define DCMAC__C8_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C8_CTL_TX_FCS_INS_ENABLE    32'h00000497
`define DCMAC__C8_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C8_CTL_TX_IGNORE_FCS    32'h00000498
`define DCMAC__C8_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C8_CTL_TX_IPG_VALUE    32'h00000499
`define DCMAC__C8_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C8_CTL_TX_SEND_IDLE    32'h0000049a
`define DCMAC__C8_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C8_CTL_TX_SEND_LFI    32'h0000049b
`define DCMAC__C8_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C8_CTL_TX_SEND_RFI    32'h0000049c
`define DCMAC__C8_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__C9_CTL_RX_CHECK_PREAMBLE    32'h0000049d
`define DCMAC__C9_CTL_RX_CHECK_PREAMBLE_SZ 40

`define DCMAC__C9_CTL_RX_CHECK_SFD    32'h0000049e
`define DCMAC__C9_CTL_RX_CHECK_SFD_SZ 40

`define DCMAC__C9_CTL_RX_DELETE_FCS    32'h0000049f
`define DCMAC__C9_CTL_RX_DELETE_FCS_SZ 40

`define DCMAC__C9_CTL_RX_IGNORE_FCS    32'h000004a0
`define DCMAC__C9_CTL_RX_IGNORE_FCS_SZ 40

`define DCMAC__C9_CTL_RX_IGNORE_INRANGE    32'h000004a1
`define DCMAC__C9_CTL_RX_IGNORE_INRANGE_SZ 40

`define DCMAC__C9_CTL_RX_IS_CLAUSE_49    32'h000004a2
`define DCMAC__C9_CTL_RX_IS_CLAUSE_49_SZ 40

`define DCMAC__C9_CTL_RX_MAX_PACKET_LEN    32'h000004a3
`define DCMAC__C9_CTL_RX_MAX_PACKET_LEN_SZ 14

`define DCMAC__C9_CTL_RX_PROCESS_LFI    32'h000004a4
`define DCMAC__C9_CTL_RX_PROCESS_LFI_SZ 40

`define DCMAC__C9_CTL_TX_CORRUPT_FCS_ON_ERR    32'h000004a5
`define DCMAC__C9_CTL_TX_CORRUPT_FCS_ON_ERR_SZ 2

`define DCMAC__C9_CTL_TX_CUSTOM_PREAMBLE_ENABLE    32'h000004a6
`define DCMAC__C9_CTL_TX_CUSTOM_PREAMBLE_ENABLE_SZ 40

`define DCMAC__C9_CTL_TX_FCS_INS_ENABLE    32'h000004a7
`define DCMAC__C9_CTL_TX_FCS_INS_ENABLE_SZ 40

`define DCMAC__C9_CTL_TX_IGNORE_FCS    32'h000004a8
`define DCMAC__C9_CTL_TX_IGNORE_FCS_SZ 40

`define DCMAC__C9_CTL_TX_IPG_VALUE    32'h000004a9
`define DCMAC__C9_CTL_TX_IPG_VALUE_SZ 4

`define DCMAC__C9_CTL_TX_SEND_IDLE    32'h000004aa
`define DCMAC__C9_CTL_TX_SEND_IDLE_SZ 40

`define DCMAC__C9_CTL_TX_SEND_LFI    32'h000004ab
`define DCMAC__C9_CTL_TX_SEND_LFI_SZ 40

`define DCMAC__C9_CTL_TX_SEND_RFI    32'h000004ac
`define DCMAC__C9_CTL_TX_SEND_RFI_SZ 40

`define DCMAC__CTL_AXI_AF_THRESH_OVERRIDE    32'h000004ad
`define DCMAC__CTL_AXI_AF_THRESH_OVERRIDE_SZ 4

`define DCMAC__CTL_MEM_CTRL    32'h000004ae
`define DCMAC__CTL_MEM_CTRL_SZ 10

`define DCMAC__CTL_MEM_DISABLE_RX_AXI_CLK    32'h000004af
`define DCMAC__CTL_MEM_DISABLE_RX_AXI_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_RX_CORE_CLK    32'h000004b0
`define DCMAC__CTL_MEM_DISABLE_RX_CORE_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_RX_FLEXIF_CLK    32'h000004b1
`define DCMAC__CTL_MEM_DISABLE_RX_FLEXIF_CLK_SZ 6

`define DCMAC__CTL_MEM_DISABLE_RX_MACIF_CLK    32'h000004b2
`define DCMAC__CTL_MEM_DISABLE_RX_MACIF_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_RX_PCS_ALIGN_BUFFER    32'h000004b3
`define DCMAC__CTL_MEM_DISABLE_RX_PCS_ALIGN_BUFFER_SZ 6

`define DCMAC__CTL_MEM_DISABLE_RX_PCS_CPCS    32'h000004b4
`define DCMAC__CTL_MEM_DISABLE_RX_PCS_CPCS_SZ 6

`define DCMAC__CTL_MEM_DISABLE_RX_PCS_DECODER    32'h000004b5
`define DCMAC__CTL_MEM_DISABLE_RX_PCS_DECODER_SZ 40

`define DCMAC__CTL_MEM_DISABLE_RX_SERDES_CLK    32'h000004b6
`define DCMAC__CTL_MEM_DISABLE_RX_SERDES_CLK_SZ 6

`define DCMAC__CTL_MEM_DISABLE_TX_AXI_CLK    32'h000004b7
`define DCMAC__CTL_MEM_DISABLE_TX_AXI_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_TX_CORE_CLK    32'h000004b8
`define DCMAC__CTL_MEM_DISABLE_TX_CORE_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_TX_FLEXIF_CLK    32'h000004b9
`define DCMAC__CTL_MEM_DISABLE_TX_FLEXIF_CLK_SZ 6

`define DCMAC__CTL_MEM_DISABLE_TX_MACIF_CLK    32'h000004ba
`define DCMAC__CTL_MEM_DISABLE_TX_MACIF_CLK_SZ 40

`define DCMAC__CTL_MEM_DISABLE_TX_PCS_CPCS    32'h000004bb
`define DCMAC__CTL_MEM_DISABLE_TX_PCS_CPCS_SZ 6

`define DCMAC__CTL_MEM_DISABLE_TX_PCS_ENCODER    32'h000004bc
`define DCMAC__CTL_MEM_DISABLE_TX_PCS_ENCODER_SZ 40

`define DCMAC__CTL_MEM_DISABLE_TX_SERDES_CLK    32'h000004bd
`define DCMAC__CTL_MEM_DISABLE_TX_SERDES_CLK_SZ 6

`define DCMAC__CTL_MEM_DISABLE_TX_TS2PHY    32'h000004be
`define DCMAC__CTL_MEM_DISABLE_TX_TS2PHY_SZ 40

`define DCMAC__CTL_REVISION    32'h000004bf
`define DCMAC__CTL_REVISION_SZ 32

`define DCMAC__CTL_RSVD0    32'h000004c0
`define DCMAC__CTL_RSVD0_SZ 32

`define DCMAC__CTL_RSVD1    32'h000004c1
`define DCMAC__CTL_RSVD1_SZ 32

`define DCMAC__CTL_RSVD2    32'h000004c2
`define DCMAC__CTL_RSVD2_SZ 32

`define DCMAC__CTL_RSVD3    32'h000004c3
`define DCMAC__CTL_RSVD3_SZ 32

`define DCMAC__CTL_RSVD4    32'h000004c4
`define DCMAC__CTL_RSVD4_SZ 32

`define DCMAC__CTL_RSVD5    32'h000004c5
`define DCMAC__CTL_RSVD5_SZ 32

`define DCMAC__CTL_RSVD6    32'h000004c6
`define DCMAC__CTL_RSVD6_SZ 32

`define DCMAC__CTL_RSVD7    32'h000004c7
`define DCMAC__CTL_RSVD7_SZ 32

`define DCMAC__CTL_RX_ALL_CH_TICK_REG_MODE_SEL    32'h000004c8
`define DCMAC__CTL_RX_ALL_CH_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__CTL_RX_AXIS_CFG    32'h000004c9
`define DCMAC__CTL_RX_AXIS_CFG_SZ 40

`define DCMAC__CTL_RX_ECC_ERR_CLEAR    32'h000004ca
`define DCMAC__CTL_RX_ECC_ERR_CLEAR_SZ 1

`define DCMAC__CTL_RX_FEC_CK_UNIQUE_FLIP    32'h000004cb
`define DCMAC__CTL_RX_FEC_CK_UNIQUE_FLIP_SZ 40

`define DCMAC__CTL_RX_FEC_ERRIND_MODE    32'h000004cc
`define DCMAC__CTL_RX_FEC_ERRIND_MODE_SZ 40

`define DCMAC__CTL_RX_INDEPENDENT_TSMAC_AND_PHY_MODE    32'h000004cd
`define DCMAC__CTL_RX_INDEPENDENT_TSMAC_AND_PHY_MODE_SZ 40

`define DCMAC__CTL_RX_MAC_DEBUG_SELECT    32'h000004ce
`define DCMAC__CTL_RX_MAC_DEBUG_SELECT_SZ 4

`define DCMAC__CTL_RX_PCS_ACTIVE_PORTS    32'h000004cf
`define DCMAC__CTL_RX_PCS_ACTIVE_PORTS_SZ 3

`define DCMAC__CTL_RX_PHY_DEBUG_SELECT    32'h000004d0
`define DCMAC__CTL_RX_PHY_DEBUG_SELECT_SZ 5

`define DCMAC__CTL_TEST_MODE_MEMCEL    32'h000004d1
`define DCMAC__CTL_TEST_MODE_MEMCEL_SZ 4

`define DCMAC__CTL_TX_ALL_CH_TICK_REG_MODE_SEL    32'h000004d2
`define DCMAC__CTL_TX_ALL_CH_TICK_REG_MODE_SEL_SZ 40

`define DCMAC__CTL_TX_AXIS_CFG    32'h000004d3
`define DCMAC__CTL_TX_AXIS_CFG_SZ 40

`define DCMAC__CTL_TX_ECC_ERR_CLEAR    32'h000004d4
`define DCMAC__CTL_TX_ECC_ERR_CLEAR_SZ 1

`define DCMAC__CTL_TX_ECC_ERR_COUNT_TICK    32'h000004d5
`define DCMAC__CTL_TX_ECC_ERR_COUNT_TICK_SZ 1

`define DCMAC__CTL_TX_FEC_CK_UNIQUE_FLIP    32'h000004d6
`define DCMAC__CTL_TX_FEC_CK_UNIQUE_FLIP_SZ 40

`define DCMAC__CTL_TX_INDEPENDENT_TSMAC_AND_PHY_MODE    32'h000004d7
`define DCMAC__CTL_TX_INDEPENDENT_TSMAC_AND_PHY_MODE_SZ 40

`define DCMAC__CTL_TX_MAC_DEBUG_SELECT    32'h000004d8
`define DCMAC__CTL_TX_MAC_DEBUG_SELECT_SZ 4

`define DCMAC__CTL_TX_PCS_ACTIVE_PORTS    32'h000004d9
`define DCMAC__CTL_TX_PCS_ACTIVE_PORTS_SZ 3

`define DCMAC__CTL_TX_PHY_DEBUG_SELECT    32'h000004da
`define DCMAC__CTL_TX_PHY_DEBUG_SELECT_SZ 4

`define DCMAC__LANE_CONNECTIVITY    32'h000004db
`define DCMAC__LANE_CONNECTIVITY_SZ 32

`define DCMAC__MAC_ACTIVITY_FACTOR    32'h000004dc
`define DCMAC__MAC_ACTIVITY_FACTOR_SZ 64

`define DCMAC__NUM_100G_FEC_NOPCS_PORTS    32'h000004dd
`define DCMAC__NUM_100G_FEC_NOPCS_PORTS_SZ 3

`define DCMAC__NUM_100G_PCS_NOFEC_PORTS    32'h000004de
`define DCMAC__NUM_100G_PCS_NOFEC_PORTS_SZ 3

`define DCMAC__NUM_100G_PCS_WITH_FEC_PORTS    32'h000004df
`define DCMAC__NUM_100G_PCS_WITH_FEC_PORTS_SZ 3

`define DCMAC__NUM_200G_PORTS    32'h000004e0
`define DCMAC__NUM_200G_PORTS_SZ 2

`define DCMAC__NUM_400G_PORTS    32'h000004e1
`define DCMAC__NUM_400G_PORTS_SZ 1

`define DCMAC__NUM_50G_FEC_NOPCS_PORTS    32'h000004e2
`define DCMAC__NUM_50G_FEC_NOPCS_PORTS_SZ 4

`define DCMAC__RXMAC_ACTIVE    32'h000004e3
`define DCMAC__RXMAC_ACTIVE_SZ 1

`define DCMAC__SIM_VERSION    32'h000004e4
`define DCMAC__SIM_VERSION_SZ 4

`define DCMAC__TXMAC_ACTIVE    32'h000004e5
`define DCMAC__TXMAC_ACTIVE_SZ 1

`endif  // B_DCMAC_DEFINES_VH