`include "B_HNICX_defines.vh"

reg [`HNICX_DATA_SZ-1:0] ATTR [0:`HNICX_ADDR_N-1];
reg [`HNICX__HNICX_DATA_RATE_SZ:1] HNICX_DATA_RATE_REG = HNICX_DATA_RATE;
reg [`HNICX__HNICX_DPU_MODE_CRYPTO_OPTIONS_SZ:1] HNICX_DPU_MODE_CRYPTO_OPTIONS_REG = HNICX_DPU_MODE_CRYPTO_OPTIONS;
reg [`HNICX__HNICX_PACKET_SIZE_SZ-1:0] HNICX_PACKET_SIZE_REG = HNICX_PACKET_SIZE;
reg [`HNICX__SIM_AES_EN_SZ:1] SIM_AES_EN_REG = SIM_AES_EN;
reg [`HNICX__SIM_CM_EN_SZ:1] SIM_CM_EN_REG = SIM_CM_EN;
reg [`HNICX__SIM_VERSION_SZ-1:0] SIM_VERSION_REG = SIM_VERSION;

initial begin
  ATTR[`HNICX__HNICX_DATA_RATE] = HNICX_DATA_RATE;
  ATTR[`HNICX__HNICX_DPU_MODE_CRYPTO_OPTIONS] = HNICX_DPU_MODE_CRYPTO_OPTIONS;
  ATTR[`HNICX__HNICX_PACKET_SIZE] = HNICX_PACKET_SIZE;
  ATTR[`HNICX__SIM_AES_EN] = SIM_AES_EN;
  ATTR[`HNICX__SIM_CM_EN] = SIM_CM_EN;
  ATTR[`HNICX__SIM_VERSION] = SIM_VERSION;
end

always @(trig_attr) begin
  HNICX_DATA_RATE_REG = ATTR[`HNICX__HNICX_DATA_RATE];
  HNICX_DPU_MODE_CRYPTO_OPTIONS_REG = ATTR[`HNICX__HNICX_DPU_MODE_CRYPTO_OPTIONS];
  HNICX_PACKET_SIZE_REG = ATTR[`HNICX__HNICX_PACKET_SIZE];
  SIM_AES_EN_REG = ATTR[`HNICX__SIM_AES_EN];
  SIM_CM_EN_REG = ATTR[`HNICX__SIM_CM_EN];
  SIM_VERSION_REG = ATTR[`HNICX__SIM_VERSION];
end

// procedures to override, read attribute values

task write_attr;
  input  [`HNICX_ADDR_SZ-1:0] addr;
  input  [`HNICX_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`HNICX_DATA_SZ-1:0] read_attr;
  input  [`HNICX_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
