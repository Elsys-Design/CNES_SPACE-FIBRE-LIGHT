// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_OUTPUT_DEFINES_VH
`else
`define B_DSP_OUTPUT_DEFINES_VH

// Look-up table parameters
//

`define DSP_OUTPUT_ADDR_N  10
`define DSP_OUTPUT_ADDR_SZ 32
`define DSP_OUTPUT_DATA_SZ 120

// Attribute addresses
//

`define DSP_OUTPUT__AUTORESET_PATDET    32'h00000000
`define DSP_OUTPUT__AUTORESET_PATDET_SZ 120

`define DSP_OUTPUT__AUTORESET_PRIORITY    32'h00000001
`define DSP_OUTPUT__AUTORESET_PRIORITY_SZ 40

`define DSP_OUTPUT__IS_CLK_INVERTED    32'h00000002
`define DSP_OUTPUT__IS_CLK_INVERTED_SZ 1

`define DSP_OUTPUT__IS_RSTP_INVERTED    32'h00000003
`define DSP_OUTPUT__IS_RSTP_INVERTED_SZ 1

`define DSP_OUTPUT__MASK    32'h00000004
`define DSP_OUTPUT__MASK_SZ 48

`define DSP_OUTPUT__PATTERN    32'h00000005
`define DSP_OUTPUT__PATTERN_SZ 48

`define DSP_OUTPUT__PREG    32'h00000006
`define DSP_OUTPUT__PREG_SZ 32

`define DSP_OUTPUT__SEL_MASK    32'h00000007
`define DSP_OUTPUT__SEL_MASK_SZ 112

`define DSP_OUTPUT__SEL_PATTERN    32'h00000008
`define DSP_OUTPUT__SEL_PATTERN_SZ 56

`define DSP_OUTPUT__USE_PATTERN_DETECT    32'h00000009
`define DSP_OUTPUT__USE_PATTERN_DETECT_SZ 72

`endif  // B_DSP_OUTPUT_DEFINES_VH