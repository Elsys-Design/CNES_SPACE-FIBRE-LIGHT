-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation data : 03/09/2024
--
-- Description :
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
   use phy_plus_lane_lib.pkg_phy_plus_lane.all;

entity rx_sync_fsm is
   port(
      CLK_SYS                              : in  std_logic;                       --! MAIN CLOCK
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP
      -- FROM Data-link layer
      LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer.
      -- TO lane_ctrl_word_detection
      DATA_RX_TO_LCWD                  : out std_logic_vector(31 downto 00);  --! 32-bit data to lane_ctrl_word_detect
      VALID_K_CHARAC_TO_LCWD            : out std_logic_vector(03 downto 00);  --! 4-bit valid K character flags to lane_ctrl_word_detect
      DATA_RDY_TO_LCWD                 : out std_logic;                       --! Data valid flag to lane_ctrl_word_detect
      -- FROM MANUFACTURER IP
      DATA_RX_FROM_IP                  : in  std_logic_vector(31 downto 00);  --! 32-bit data from GTY IP
      VALID_K_CHARAC_FROM_IP            : in  std_logic_vector(03 downto 00);  --! 4-bit valid K character flags from GTY IP
      DATA_RDY_FROM_IP                 : in  std_logic;                       --! Data valid flag from GTY IP
      INVALID_CHAR_FROM_IP             : in  std_logic_vector(03 downto 00);  --! Invalid character flags from GTY IP
      DISPARITY_ERR_FROM_IP            : in  std_logic_vector(03 downto 00);  --! Disparity error flags from GTY IP
      RX_WORD_REALIGN_FROM_IP          : in  std_logic;                       --! RX word realign from GTY IP
      COMMA_DET_FROM_IP                : in  std_logic;                       --! Flag indicates that a comma is detected on the word receive
      -- PARAMETERS
      LANE_RESET                       : in  std_logic                        --! Asserts or de-asserts LaneReset for the lane
   );
end rx_sync_fsm;

architecture rtl of rx_sync_fsm is

----------------------------- Declaration signals -----------------------------
-- Receiver synchronisation FSM transition conditions process
   -- Type
type rx_sync_fsm_type is (
   LOST_SYNC_ST,                                                           --! IDLE state of the FSM
   CHECK_SYNC_ST,                                                          --! Checking data to validate synchronisation state
   READY_ST                                                                --! Synchronisation ok state
   );
   -- Signals
signal current_state                : rx_sync_fsm_type;                    --! Current state of the Lane Initialisation FSM
signal comma_det_from_ip_r          : std_logic;                           --! COMMA_DET_FROM_IP registered signal
signal rx_word_realign_from_ip_r    : std_logic;                           --! word realignement flag registered
signal rx_word_realign_from_ip_rr    : std_logic;                           --! word realignement flag registered bis
signal data_rx_to_lcwd_i            : std_logic_vector(31 downto 00);      --! 32-bit data send to lane_ctrl_word_detect
signal valid_k_charac_to_lcwd_i     : std_logic_vector(03 downto 00);      --! 4-bit valid K character flags to lane_ctrl_word_detect
signal data_rdy_to_lcwd_i           : std_logic;                           --! Data valid flag to lane_ctrl_word_detect
signal err_word_cnt                 : unsigned(02 downto 00);              --! RXERR control word counter
signal err_word_x5                  : std_logic;                           --! Flag indicates that err_word_cnt reaches 5
signal valid_symb                   : std_logic;                           --! Flag indicates that a valid symbol is received
signal invalid_symb                 : std_logic;                           --! Flag indicates that an invalid symbol is received
signal disparity_err                : std_logic;                           --! Flag indicates that a disparity error is detected
signal test_state : std_logic_vector(1 downto 0);

begin

   -- Receiver word synchronisation FSM tansition process
   p_rx_sync_fsm_transition : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         current_state              <= LOST_SYNC_ST;
         rx_word_realign_from_ip_r  <= '0';
         rx_word_realign_from_ip_rr <= '0';
         comma_det_from_ip_r        <= '0';
         test_state <="00";
      elsif rising_edge(CLK) then
         rx_word_realign_from_ip_r  <= RX_WORD_REALIGN_FROM_IP;
         rx_word_realign_from_ip_rr <= rx_word_realign_from_ip_r;
         comma_det_from_ip_r        <= COMMA_DET_FROM_IP;

         case current_state is

            when LOST_SYNC_ST   =>  if (COMMA_DET_FROM_IP = '1' and comma_det_from_ip_r = '0')  or COMMA_DET_FROM_IP = '1' then  -- when a Comma sequence is detected
                                       current_state  <= CHECK_SYNC_ST;                            -- FSM goes to next state
                                    else                                                           -- else
                                       current_state  <= LOST_SYNC_ST;                             -- Stays in current state
                                    end if;
                                    test_state <="00";


            when CHECK_SYNC_ST  =>  if (LANE_RESET = '1' or LANE_RESET_DL = '1')  or ((rx_word_realign_from_ip_r = '1' and rx_word_realign_from_ip_rr = '0') or rx_word_realign_from_ip_r = '1') or err_word_x5 = '1' then
                                       current_state  <= LOST_SYNC_ST;
                                    elsif valid_symb = '1' then
                                       current_state  <= READY_ST;
                                    else
                                       current_state  <= CHECK_SYNC_ST;
                                    end if;
                                    test_state <="01";


            when READY_ST       =>  if (LANE_RESET = '1' or LANE_RESET_DL = '1') or ((rx_word_realign_from_ip_r = '1' and rx_word_realign_from_ip_rr = '0') or rx_word_realign_from_ip_r = '1') then
                                       current_state  <= LOST_SYNC_ST;
                                    elsif invalid_symb = '1' or disparity_err = '1' then
                                       current_state  <= CHECK_SYNC_ST;
                                    else
                                       current_state  <= READY_ST;
                                    end if;
                                    test_state <="11";

            when others          => current_state  <= LOST_SYNC_ST;

         end case;
      end if;
   end process p_rx_sync_fsm_transition;

   -- Receiver word synchronisation FSM actions on state process
   p_rx_sync_action_on_state : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         data_rx_to_lcwd_i          <= (others => '0');
         valid_k_charac_to_lcwd_i   <= (others => '0');
         data_rdy_to_lcwd_i         <= '0';
         err_word_cnt               <= (others => '0');
         err_word_x5                <= '0';
         valid_symb                 <= '0';
         invalid_symb               <= '0';
         disparity_err              <= '0';

      elsif rising_edge(CLK) then

         if current_state = LOST_SYNC_ST then

            err_word_cnt               <= (others => '0');           -- reset counter
            err_word_x5                <= '0';                       -- De-asserts flag
            data_rx_to_lcwd_i          <= C_RXERR_WORD;              -- Replace data receive by RX_ERR control word
            valid_k_charac_to_lcwd_i   <= x"1";                      -- All word symbol are K character
            data_rdy_to_lcwd_i         <= '1';                       -- Asserts handshake


         elsif current_state = CHECK_SYNC_ST then

            invalid_symb      <= '0';                                -- De-asserts flag
            disparity_err     <= '0';                                -- De-asserts flag

            if DATA_RDY_FROM_IP = '1' then                           -- when a data is receive from MANUFACTURER IP

               data_rx_to_lcwd_i          <= DATA_RX_FROM_IP;        -- Data from IP is send to lane_ctrl_word_detection
               valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_FROM_IP;  -- Valid K character from IP is send to lane_ctrl_word_detection
               data_rdy_to_lcwd_i         <= '1';                    -- Asserts handshake

               if INVALID_CHAR_FROM_IP /= x"0" or DISPARITY_ERR_FROM_IP /= x"0" then   -- When only one Symbol of the 32-bit word is an invalid character or disparity error
                  data_rx_to_lcwd_i          <= C_RXERR_WORD;              -- Replace data receive by RX_ERR control word
                  valid_k_charac_to_lcwd_i   <= x"1";                      -- All word symbol are K character
                  if err_word_cnt >= C_SYMB_X5 then                                    -- and 5 characters cointaining an error has been received consecultively
                     err_word_x5   <= '1';                                             -- Asserts flag
                  elsif err_word_cnt < C_SYMB_X5 then                                  -- else
                     err_word_cnt  <= err_word_cnt + 1;                                -- increment counter
                     err_word_x5   <= '0';                                             -- De-asserts flag
                  end if;
               else
                  valid_symb    <= '1';                                                -- Asserts flag
                  err_word_cnt  <= (others => '0');                                    -- reset error flag and counter
                  err_word_x5   <= '0';
               end if;

            else
               data_rx_to_lcwd_i          <= (others => '0');        -- Data from IP is reseted
               valid_k_charac_to_lcwd_i   <= (others => '0');        -- Valid K character is reseted
               data_rdy_to_lcwd_i         <= '0';                    -- De-asserts handshake
            end if;

         elsif current_state = READY_ST then

            err_word_cnt         <= (others => '0');                 -- reset counter
            valid_symb           <= '0';                             -- De-asserts flag
            if DATA_RDY_FROM_IP = '1' then                           -- when a data is receive from MANUFACTURER IP

               data_rx_to_lcwd_i          <= DATA_RX_FROM_IP;        -- Data from IP is send to lane_ctrl_word_detection
               valid_k_charac_to_lcwd_i   <= VALID_K_CHARAC_FROM_IP;  -- Valid K character from IP is send to lane_ctrl_word_detection
               data_rdy_to_lcwd_i         <= '1';                    -- Asserts handshake

               if INVALID_CHAR_FROM_IP /= x"0" then                     -- When only one Symbol of the 32-bit word is an invalid character
                  invalid_symb      <= '1';                             -- Asserts flag
                  data_rx_to_lcwd_i          <= C_RXERR_WORD;              -- Replace data receive by RX_ERR control word
                  valid_k_charac_to_lcwd_i   <= x"1";                      -- All word symbol are K character
               else                                                     -- else
                  invalid_symb      <= '0';                             -- De-asserts flag
               end if;

               if DISPARITY_ERR_FROM_IP /= x"0" then                    -- When only one Symbol of the 32-bit word is an disparity error
                  disparity_err     <= '1';                             -- Asserts flag
                  data_rx_to_lcwd_i          <= C_RXERR_WORD;              -- Replace data receive by RX_ERR control word
                  valid_k_charac_to_lcwd_i   <= x"1";                      -- All word symbol are K character
               else                                                     -- else
                  disparity_err     <= '0';                             -- De-asserts flag
               end if;
            end if;
         end if;
      end if;
   end process p_rx_sync_action_on_state;


-- Outputs
DATA_RX_TO_LCWD         <= data_rx_to_lcwd_i;
VALID_K_CHARAC_TO_LCWD   <= valid_k_charac_to_lcwd_i;
DATA_RDY_TO_LCWD        <= data_rdy_to_lcwd_i;

end architecture rtl;
