`include "B_HBM_SNGLBLI_INTF_AXI_defines.vh"

reg [`HBM_SNGLBLI_INTF_AXI_DATA_SZ-1:0] ATTR [0:`HBM_SNGLBLI_INTF_AXI_ADDR_N-1];
reg [`HBM_SNGLBLI_INTF_AXI__CLK_SEL_SZ:1] CLK_SEL_REG = CLK_SEL;
reg [`HBM_SNGLBLI_INTF_AXI__DATARATE_SZ-1:0] DATARATE_REG = DATARATE;
reg IS_ACLK_INVERTED_REG = IS_ACLK_INVERTED;
reg IS_ARESET_N_INVERTED_REG = IS_ARESET_N_INVERTED;
reg [`HBM_SNGLBLI_INTF_AXI__MC_ENABLE_SZ:1] MC_ENABLE_REG = MC_ENABLE;
reg [`HBM_SNGLBLI_INTF_AXI__PAGEHIT_PERCENT_SZ-1:0] PAGEHIT_PERCENT_REG = PAGEHIT_PERCENT;
reg [`HBM_SNGLBLI_INTF_AXI__PHY_ENABLE_SZ:1] PHY_ENABLE_REG = PHY_ENABLE;
reg [`HBM_SNGLBLI_INTF_AXI__READ_PERCENT_SZ-1:0] READ_PERCENT_REG = READ_PERCENT;
reg [`HBM_SNGLBLI_INTF_AXI__SWITCH_ENABLE_SZ:1] SWITCH_ENABLE_REG = SWITCH_ENABLE;
reg [`HBM_SNGLBLI_INTF_AXI__WRITE_PERCENT_SZ-1:0] WRITE_PERCENT_REG = WRITE_PERCENT;

initial begin
  ATTR[`HBM_SNGLBLI_INTF_AXI__CLK_SEL] = CLK_SEL;
  ATTR[`HBM_SNGLBLI_INTF_AXI__DATARATE] = DATARATE;
  ATTR[`HBM_SNGLBLI_INTF_AXI__IS_ACLK_INVERTED] = IS_ACLK_INVERTED;
  ATTR[`HBM_SNGLBLI_INTF_AXI__IS_ARESET_N_INVERTED] = IS_ARESET_N_INVERTED;
  ATTR[`HBM_SNGLBLI_INTF_AXI__MC_ENABLE] = MC_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_AXI__PAGEHIT_PERCENT] = PAGEHIT_PERCENT;
  ATTR[`HBM_SNGLBLI_INTF_AXI__PHY_ENABLE] = PHY_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_AXI__READ_PERCENT] = READ_PERCENT;
  ATTR[`HBM_SNGLBLI_INTF_AXI__SWITCH_ENABLE] = SWITCH_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_AXI__WRITE_PERCENT] = WRITE_PERCENT;
end

always @(trig_attr) begin
  CLK_SEL_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__CLK_SEL];
  DATARATE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__DATARATE];
  IS_ACLK_INVERTED_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__IS_ACLK_INVERTED];
  IS_ARESET_N_INVERTED_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__IS_ARESET_N_INVERTED];
  MC_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__MC_ENABLE];
  PAGEHIT_PERCENT_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__PAGEHIT_PERCENT];
  PHY_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__PHY_ENABLE];
  READ_PERCENT_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__READ_PERCENT];
  SWITCH_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__SWITCH_ENABLE];
  WRITE_PERCENT_REG = ATTR[`HBM_SNGLBLI_INTF_AXI__WRITE_PERCENT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`HBM_SNGLBLI_INTF_AXI_ADDR_SZ-1:0] addr;
  input  [`HBM_SNGLBLI_INTF_AXI_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`HBM_SNGLBLI_INTF_AXI_DATA_SZ-1:0] read_attr;
  input  [`HBM_SNGLBLI_INTF_AXI_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
