------------------------------------------------------------------------
--
-- Copyright 1996 by IEEE. All rights reserved.
--
-- This source file is an essential part of IEEE Std 1076.2-1996, IEEE Standard
-- VHDL Mathematical Packages. This source file may not be copied, sold, or
-- included with software that is sold without written permission from the IEEE
-- Standards Department. This source file may be used to implement this standard
-- and may be distributed in compiled form in any manner so long as the
-- compiled form does not allow direct decompilation of the original source file.
-- This source file may be copied for individual use between licensed users.
-- This source file is provided on an AS IS basis. The IEEE disclaims ANY
-- WARRANTY EXPRESS OR IMPLIED INCLUDING ANY WARRANTY OF MERCHANTABILITY
-- AND FITNESS FOR USE FOR A PARTICULAR PURPOSE. The user of the source
-- file shall indemnify and hold IEEE harmless from any damages or liability
-- arising out of the use thereof.
--
-- Title:       Standard VHDL Mathematical Packages (IEEE Std 1076.2-1996,
--              MATH_REAL)
--
-- Library:     This package shall be compiled into a library
--              symbolically named IEEE.
--
-- Developers:  IEEE DASC VHDL Mathematical Packages Working Group
--
-- Purpose:     This package defines a standard for designers to use in
--              describing VHDL models that make use of common REAL constants
--              and common REAL elementary mathematical functions.
--
-- Limitation:  The values generated by the functions in this package may
--              vary from platform to platform, and the precision of results
--              is only guaranteed to be the minimum required by IEEE Std 1076-
--              1993.
--
-- Notes:
--              No declarations or definitions shall be included in, or
--              excluded from, this package.
--              The "package declaration" defines the types, subtypes, and
--              declarations of MATH_REAL.
--              The standard mathematical definition and conventional meaning
--              of the mathematical functions that are part of this standard
--              represent the formal semantics of the implementation of the
--              MATH_REAL package declaration.  The purpose of the MATH_REAL
--              package body is to provide a guideline for implementations to
--              verify their implementation of MATH_REAL.  Tool developers may
--              choose to implement the package body in the most efficient
--              manner available to them.
--
-- -----------------------------------------------------------------------------
-- Version    : 1.5
-- Date       : 24 July 1996
-- -----------------------------------------------------------------------------

package math_real is
    constant CopyRightNotice: string
      := "Copyright 1996 IEEE. All rights reserved.";

    -- Constant Definitions

    constant MATH_E             : real := 2.71828_18284_59045_23536; -- Value of e
    constant MATH_1_OVER_E      : real := 0.36787_94411_71442_32160; -- Value of 1/e
    constant MATH_PI            : real := 3.14159_26535_89793_23846; -- Value of pi
    constant MATH_2_PI          : real := 6.28318_53071_79586_47693; -- Value of 2*pi
    constant MATH_1_OVER_PI     : real := 0.31830_98861_83790_67154; -- Value of 1/pi
    constant MATH_PI_OVER_2     : real := 1.57079_63267_94896_61923; -- Value of pi/2
    constant MATH_PI_OVER_3     : real := 1.04719_75511_96597_74615; -- Value of pi/3
    constant MATH_PI_OVER_4     : real := 0.78539_81633_97448_30962; -- Value of pi/4
    constant MATH_3_PI_OVER_2   : real := 4.71238_89803_84689_85769; -- Value 3*pi/2
    constant MATH_LOG_OF_2      : real := 0.69314_71805_59945_30942; -- Natural log of 2
    constant MATH_LOG_OF_10     : real := 2.30258_50929_94045_68402; -- Natural log of 10
    constant MATH_LOG2_OF_E     : real := 1.44269_50408_88963_4074; -- Log base 2 of e
    constant MATH_LOG10_OF_E    : real := 0.43429_44819_03251_82765; -- Log base 10 of e
    constant MATH_SQRT_2        : real := 1.41421_35623_73095_04880; -- square root of 2
    constant MATH_1_OVER_SQRT_2 : real := 0.70710_67811_86547_52440; -- square root of 1/2
    constant MATH_SQRT_PI       : real := 1.77245_38509_05516_02730; -- square root of pi
    constant MATH_DEG_TO_RAD    : real := 0.01745_32925_19943_29577; -- Conversion factor from degree to radian
    constant MATH_RAD_TO_DEG    : real := 57.29577_95130_82320_87680; -- Conversion factor from radian to degree


    -- Function Declarations

    --```
    -- Purpose:
    --         Returns 1.0 if x > 0.0; 0.0 if x = 0.0; -1.0 if x < 0.0
    -- Special values:
    --         None
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         abs(sign(x)) <= 1.0
    -- Notes:
    --         None
    --```
    function sign (x: in real ) return real;

    --```
    -- Purpose:
    --         Returns smallest integer value (as real) not less than x
    -- Special values:
    --         None
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         ceil(x) is mathematically unbounded
    -- Notes:
    --         a) Implementations have to support at least the domain
    --                abs(x) < real(integer'high)
    --```
    function ceil (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns largest integer value (as real) not greater than x
    -- Special values:
    --         floor(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         floor(x) is mathematically unbounded
    -- Notes:
    --         a) Implementations have to support at least the domain
    --                abs(x) < real(integer'high)
    --```
    function floor (x : in real ) return real;

    --```
    -- Purpose:
    --         Rounds x to the nearest integer value (as real). if x is
    --         halfway between two integers, rounding is away from 0.0
    -- Special values:
    --         round(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         round(x) is mathematically unbounded
    -- Notes:
    --         a) Implementations have to support at least the domain
    --                abs(x) < real(integer'high)
    --```
    function round (x : in real ) return real;

    --```
    -- Purpose:
    --         Truncates x towards 0.0 and returns truncated value
    -- Special values:
    --         trunc(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         trunc(x) is mathematically unbounded
    -- Notes:
    --         a) Implementations have to support at least the domain
    --                abs(x) < real(integer'high)
    --```
    function trunc (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns floating point modulus of x/y, with the same sign as
    --         y, and absolute value less than the absolute value of y, and
    --         for some integer value n the result satisfies the relation
    --         x = y*n + mod(x,y)
    -- Special values:
    --         None
    -- Domain:
    --         x in real; y in real and y /= 0.0
    -- Error conditions:
    --         Error if y = 0.0
    -- Range:
    --         abs(mod(x,y)) < abs(y)
    -- Notes:
    --         None
    --```
    function "mod" (x, y: in real ) return real;

    --```
    -- Purpose:
    --         Returns the algebraically larger of x and y
    -- Special values:
    --         realmax(x,y) = x when x = y
    -- Domain:
    --         x in real; y in real
    -- Error conditions:
    --         None
    -- Range:
    --         realmax(x,y) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function realmax (x, y : in real ) return real;

    --```
    -- Purpose:
    --         Returns the algebraically smaller of x and y
    -- Special values:
    --         realmin(x,y) = x when x = y
    -- Domain:
    --         x in real; y in real
    -- Error conditions:
    --         None
    -- Range:
    --         realmin(x,y) is mathematically unbounded
    -- Notes:
    --         None
    --```
    function realmin (x, y : in real ) return real;

    --```
    -- Purpose:
    --         Returns, in x, a pseudo-random number with uniform
    --         distribution in the open interval (0.0, 1.0).
    -- Special values:
    --         None
    -- Domain:
    --         1 <= SEED1 <= 2147483562; 1 <= SEED2 <= 2147483398
    -- Error conditions:
    --         Error if SEED1 or SEED2 outside of valid domain
    -- Range:
    --         0.0 < x < 1.0
    -- Notes:
    --         a) The semantics for this function are described by the
    --            algorithm published by Pierre L'Ecuyer in "Communications
    --            of the ACM," vol. 31, no. 6, June 1988, pp. 742-774.
    --            The algorithm is based on the combination of two
    --            multiplicative linear congruential generators for 32-bit
    --            platforms.
    --
    --         b) Before the first call to UNIFORM, the seed values
    --            (SEED1, SEED2) have to be initialized to values in the range
    --            [1, 2147483562] and [1, 2147483398] respectively.  The
    --            seed values are modified after each call to UNIFORM.
    --
    --         c) This random number generator is portable for 32-bit
    --            computers, and it has a period of ~2.30584*(10**18) for each
    --            set of seed values.
    --
    --         d) For information on spectral tests for the algorithm, refer
    --            to the L'Ecuyer article.
    --```
    procedure uniform(variable seed1,seed2:inout positive; variable x:out real);

    --```
    -- Purpose:
    --         Returns square root of x
    -- Special values:
    --         sqrt(0.0) = 0.0
    --         sqrt(1.0) = 1.0
    -- Domain:
    --         x >= 0.0
    -- Error conditions:
    --         Error if X < 0.0
    -- Range:
    --         sqrt(x) >= 0.0
    -- Notes:
    --         a) The upper bound of the reachable range of sqrt is
    --            approximately given by:
    --                sqrt(x) <= sqrt(real'high)
    --```
    function sqrt (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns cube root of x
    -- Special values:
    --         cbrt(0.0) = 0.0
    --         cbrt(1.0) = 1.0
    --         cbrt(-1.0) = -1.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         cbrt(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of cbrt is approximately given by:
    --                abs(cbrt(x)) <= cbrt(real'high)
    --```
    function cbrt (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns y power of x ==>  x**y
    -- Special values:
    --         x**0.0 = 1.0; x /= 0
    --         0**y = 0.0; y > 0.0
    --         x**1.0 = real(x); x >= 0
    --         1**y = 1.0
    -- Domain:
    --         x > 0
    --         x = 0 for y > 0.0
    --         x < 0 for y = 0.0
    -- Error conditions:
    --         Error if X < 0 and Y /= 0.0
    --         Error if X = 0 and Y <= 0.0
    -- Range:
    --         x**y >= 0.0
    -- Notes:
    --         a) The upper bound of the reachable range for "**" is
    --            approximately given by:
    --                x**y <= real'high
    --```
    function "**" (x : in integer; y : in real) return real;

    --```
    -- Purpose:
    --         Returns y power of x ==>  x**y
    -- Special values:
    --         x**0.0 = 1.0; x /= 0.0
    --         0.0**y = 0.0; y > 0.0
    --         x**1.0 = x; x >= 0.0
    --         1.0**y = 1.0
    -- Domain:
    --         x > 0.0
    --         x = 0.0 for y > 0.0
    --         x < 0.0 for y = 0.0
    -- Error conditions:
    --         Error if x < 0.0 and y /= 0.0
    --         Error if x = 0.0 and y <= 0.0
    -- Range:
    --         x**y >= 0.0
    -- Notes:
    --         a) The upper bound of the reachable range for "**" is
    --            approximately given by:
    --                x**y <= real'high
    --```
    function "**" (x : in real; y : in real) return real;

    --```
    -- Purpose:
    --         Returns e**x; where e = math_e
    -- Special values:
    --         exp(0.0) = 1.0
    --         exp(1.0) = math_e
    --         exp(-1.0) = math_1_over_e
    --         exp(x) = 0.0 for x <= -log(real'high)
    -- Domain:
    --         x in real such that exp(x) <= real'high
    -- Error conditions:
    --         Error if x > log(real'high)
    -- Range:
    --         exp(x) >= 0.0
    -- Notes:
    --         a) The usable domain of exp is approximately given by:
    --                x <= log(real'high)
    --```
    function exp (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns natural logarithm of x
    -- Special values:
    --         log(1.0) = 0.0
    --         log(math_e) = 1.0
    -- Domain:
    --         x > 0.0
    -- Error conditions:
    --         Error if x <= 0.0
    -- Range:
    --         log(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of log is approximately given by:
    --                log(0+) <= log(x) <= log(real'high)
    --```
    function log (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns logarithm base 2 of x
    -- Special values:
    --         log2(1.0) = 0.0
    --         log2(2.0) = 1.0
    -- Domain:
    --         x > 0.0
    -- Error conditions:
    --         Error if x <= 0.0
    -- Range:
    --         log2(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of log2 is approximately given by:
    --                log2(0+) <= log2(x) <= log2(real'high)
    --```
    function log2 (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns logarithm base 10 of x
    -- Special values:
    --         log10(1.0) = 0.0
    --         log10(10.0) = 1.0
    -- Domain:
    --         x > 0.0
    -- Error conditions:
    --         Error if x <= 0.0
    -- Range:
    --         log10(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of log10 is approximately given by:
    --                Log10(0+) <= log10(x) <= log10(real'high)
    --```
    function log10 (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns logarithm base base of x
    -- Special values:
    --         log(1.0, base) = 0.0
    --         log(base, base) = 1.0
    -- Domain:
    --         x > 0.0
    --         base > 0.0
    --         base /= 1.0
    -- Error conditions:
    --         Error if x <= 0.0
    --         Error if base <= 0.0
    --         Error if base = 1.0
    -- Range:
    --         log(x, base) is mathematically unbounded
    -- Notes:
    --         a) When base > 1.0, the reachable range of log is
    --            approximately given by:
    --                log(0+, base) <= log(x, base) <= log(real'high, base)
    --         b) When 0.0 < base < 1.0, the reachable range of log is
    --            approximately given by:
    --                log(real'high, base) <= log(x, base) <= log(0+, base)
    --```
    function log (x: in real; base: in real) return real;

    --```
    -- Purpose:
    --         Returns sine of x; x in radians
    -- Special values:
    --         sin(x) = 0.0 for x = k*MATH_PI, where k is an integer
    --         sin(x) = 1.0 for x = (4*k+1)*MATH_PI_OVER_2, where k is an integer
    --         sin(x) = -1.0 for x = (4*k+3)*MATH_PI_OVER_2, where k is an integer
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         abs(sin(x)) <= 1.0
    -- Notes:
    --         a) For larger values of abs(x), degraded accuracy is allowed.
    --```
    function  sin (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns cosine of x; x in radians
    -- Special values:
    --         cos(x) = 0.0 for x = (2*k+1)*MATH_PI_OVER_2, where k is an integer
    --         cos(x) = 1.0 for x = (2*k)*MATH_PI, where k is an integer
    --         cos(x) = -1.0 for x = (2*k+1)*MATH_PI, where k is an integer
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         abs(cos(x)) <= 1.0
    -- Notes:
    --         a) For larger values of abs(x), degraded accuracy is allowed.
    --```
    function  cos ( x : in real ) return real;

    --```
    -- Purpose:
    --         Returns tangent of x; x in radians
    -- Special values:
    --         tan(x) = 0.0 for x = k*MATH_PI, where k is an integer
    -- Domain:
    --         x in real and
    --         x /= (2*k+1)*MATH_PI_OVER_2, where k is an integer
    -- Error conditions:
    --         Error if x = ((2*k+1) * MATH_PI_OVER_2), where k is an integer
    -- Range:
    --         tan(x) is mathematically unbounded
    -- Notes:
    --         a) For larger values of abs(x), degraded accuracy is allowed.
    --```
    function  tan (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns inverse sine of x
    -- Special values:
    --         arcsin(0.0) = 0.0
    --         arcsin(1.0) = MATH_PI_OVER_2
    --         arcsin(-1.0) = -MATH_PI_OVER_2
    -- Domain:
    --         abs(x) <= 1.0
    -- Error conditions:
    --         Error if abs(x) > 1.0
    -- Range:
    --         abs(arcsin(x) <= MATH_PI_OVER_2
    -- Notes:
    --         None
    --```
    function  arcsin (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns inverse cosine of x
    -- Special values:
    --         arccos(1.0) = 0.0
    --         arccos(0.0) = MATH_PI_OVER_2
    --         arccos(-1.0) = MATH_PI
    -- Domain:
    --         abs(x) <= 1.0
    -- Error conditions:
    --         Error if ABS(X) > 1.0
    -- Range:
    --         0.0 <= arccos(x) <= MATH_PI
    -- Notes:
    --         None
    --```
    function  arccos (x : in real ) return real;

    --```
    -- Purpose:
    --         Returns the value of the angle in radians of the point
    --        (1.0, Y), which is in rectangular coordinates
    -- Special values:
    --         arctan(0.0) = 0.0
    -- Domain:
    --         y in real
    -- Error conditions:
    --         None
    -- Range:
    --         abs(arctan(y)) <= MATH_PI_OVER_2
    -- Notes:
    --         None
    --```
    function  arctan (y : in real) return real;

    --```
    -- Purpose:
    --         Returns the principal value of the angle in radians of
    --         the point (X, Y), which is in rectangular coordinates
    -- Special values:
    --         arctan(0.0, x) = 0.0 if x > 0.0
    --         arctan(0.0, x) = MATH_PI if x < 0.0
    --         arctan(y, 0.0) = MATH_PI_OVER_2 if y > 0.0
    --         arctan(y, 0.0) = -MATH_PI_OVER_2 if y < 0.0
    -- Domain:
    --         y in real
    --         x in real, x /= 0.0 when y = 0.0
    -- Error conditions:
    --         Error if X = 0.0 and Y = 0.0
    -- Range:
    --         -MATH_PI < arctan(y,x) <= MATH_PI
    -- Notes:
    --         None
    --```
    function  arctan (y : in real; x : in real) return real;

    --```
    -- Purpose:
    --         Returns hyperbolic sine of x
    -- Special values:
    --         sinh(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         sinh(x) is mathematically unbounded
    -- Notes:
    --         a) The usable domain of sinh is approximately given by:
    --                abs(x) <= log(real'high)
    --```
    function sinh (x : in real) return real;

    --```
    -- Purpose:
    --         Returns hyperbolic cosine of x
    -- Special values:
    --         cosh(0.0) = 1.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         cosh(x) >= 1.0
    -- Notes:
    --         a) The usable domain of cosh is approximately given by:
    --                abs(x) <= log(real'high)
    --```
    function cosh (x : in real) return real;

    --```
    -- Purpose:
    --         Returns hyperbolic tangent of x
    -- Special values:
    --         tanh(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         abs(tanh(x)) <= 1.0
    -- Notes:
    --         None
    --```
    function tanh (x : in real) return real;

    --```
    -- Purpose:
    --         Returns inverse hyperbolic sine of x
    -- Special values:
    --         arcsinh(0.0) = 0.0
    -- Domain:
    --         x in real
    -- Error conditions:
    --         None
    -- Range:
    --         arcsinh(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of arcsinh is approximately given by:
    --                abs(arcsinh(x)) <= log(real'high)
    --```
    function arcsinh (x : in real) return real;

    --```
    -- Purpose:
    --         Returns inverse hyperbolic cosine of x
    -- Special values:
    --         arccosh(1.0) = 0.0
    -- Domain:
    --         x >= 1.0
    -- Error conditions:
    --         Error if x < 1.0
    -- Range:
    --         arccosh(x) >= 0.0
    -- Notes:
    --         a) The upper bound of the reachable range of arccosh is
    --            approximately given by:   arccosh(x) <= log(real'high)
    --```
    function arccosh (x : in real) return real;

    --```
    -- Purpose:
    --         Returns inverse hyperbolic tangent of x
    -- Special values:
    --         arctanh(0.0) = 0.0
    -- Domain:
    --         abs(x) < 1.0
    -- Error conditions:
    --         Error if abs(x) >= 1.0
    -- Range:
    --         arctanh(x) is mathematically unbounded
    -- Notes:
    --         a) The reachable range of arctanh is approximately given by:
    --                abs(arctanh(x)) < log(real'high)
    --```
    function arctanh (x : in real) return real;

end package math_real;
