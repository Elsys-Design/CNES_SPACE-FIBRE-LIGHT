// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTYP_QUAD_DEFINES_VH
`else
`define B_GTYP_QUAD_DEFINES_VH

// Look-up table parameters
//

`define GTYP_QUAD_ADDR_N  792
`define GTYP_QUAD_ADDR_SZ 32
`define GTYP_QUAD_DATA_SZ 192

// Attribute addresses
//

`define GTYP_QUAD__A_CFG0    32'h00000000
`define GTYP_QUAD__A_CFG0_SZ 32

`define GTYP_QUAD__A_CFG1    32'h00000001
`define GTYP_QUAD__A_CFG1_SZ 32

`define GTYP_QUAD__A_CFG2    32'h00000002
`define GTYP_QUAD__A_CFG2_SZ 32

`define GTYP_QUAD__A_CFG3    32'h00000003
`define GTYP_QUAD__A_CFG3_SZ 32

`define GTYP_QUAD__A_CFG4    32'h00000004
`define GTYP_QUAD__A_CFG4_SZ 32

`define GTYP_QUAD__A_CFG5    32'h00000005
`define GTYP_QUAD__A_CFG5_SZ 32

`define GTYP_QUAD__CH0_ADAPT_APT_CFG    32'h00000006
`define GTYP_QUAD__CH0_ADAPT_APT_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_CAL_CFG    32'h00000007
`define GTYP_QUAD__CH0_ADAPT_CAL_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_DFE_CFG    32'h00000008
`define GTYP_QUAD__CH0_ADAPT_DFE_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GC_CFG0    32'h00000009
`define GTYP_QUAD__CH0_ADAPT_GC_CFG0_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GC_CFG1    32'h0000000a
`define GTYP_QUAD__CH0_ADAPT_GC_CFG1_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GC_CFG2    32'h0000000b
`define GTYP_QUAD__CH0_ADAPT_GC_CFG2_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GC_CFG3    32'h0000000c
`define GTYP_QUAD__CH0_ADAPT_GC_CFG3_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GEN_CFG0    32'h0000000d
`define GTYP_QUAD__CH0_ADAPT_GEN_CFG0_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GEN_CFG1    32'h0000000e
`define GTYP_QUAD__CH0_ADAPT_GEN_CFG1_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GEN_CFG2    32'h0000000f
`define GTYP_QUAD__CH0_ADAPT_GEN_CFG2_SZ 32

`define GTYP_QUAD__CH0_ADAPT_GEN_CFG3    32'h00000010
`define GTYP_QUAD__CH0_ADAPT_GEN_CFG3_SZ 32

`define GTYP_QUAD__CH0_ADAPT_H01_CFG    32'h00000011
`define GTYP_QUAD__CH0_ADAPT_H01_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_H23_CFG    32'h00000012
`define GTYP_QUAD__CH0_ADAPT_H23_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_H45_CFG    32'h00000013
`define GTYP_QUAD__CH0_ADAPT_H45_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_H67_CFG    32'h00000014
`define GTYP_QUAD__CH0_ADAPT_H67_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_H89_CFG    32'h00000015
`define GTYP_QUAD__CH0_ADAPT_H89_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_HAB_CFG    32'h00000016
`define GTYP_QUAD__CH0_ADAPT_HAB_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_HCD_CFG    32'h00000017
`define GTYP_QUAD__CH0_ADAPT_HCD_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_HEF_CFG    32'h00000018
`define GTYP_QUAD__CH0_ADAPT_HEF_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG0    32'h00000019
`define GTYP_QUAD__CH0_ADAPT_KH_CFG0_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG1    32'h0000001a
`define GTYP_QUAD__CH0_ADAPT_KH_CFG1_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG2    32'h0000001b
`define GTYP_QUAD__CH0_ADAPT_KH_CFG2_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG3    32'h0000001c
`define GTYP_QUAD__CH0_ADAPT_KH_CFG3_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG4    32'h0000001d
`define GTYP_QUAD__CH0_ADAPT_KH_CFG4_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KH_CFG5    32'h0000001e
`define GTYP_QUAD__CH0_ADAPT_KH_CFG5_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KL_CFG0    32'h0000001f
`define GTYP_QUAD__CH0_ADAPT_KL_CFG0_SZ 32

`define GTYP_QUAD__CH0_ADAPT_KL_CFG1    32'h00000020
`define GTYP_QUAD__CH0_ADAPT_KL_CFG1_SZ 32

`define GTYP_QUAD__CH0_ADAPT_LCK_CFG0    32'h00000021
`define GTYP_QUAD__CH0_ADAPT_LCK_CFG0_SZ 32

`define GTYP_QUAD__CH0_ADAPT_LCK_CFG1    32'h00000022
`define GTYP_QUAD__CH0_ADAPT_LCK_CFG1_SZ 32

`define GTYP_QUAD__CH0_ADAPT_LCK_CFG2    32'h00000023
`define GTYP_QUAD__CH0_ADAPT_LCK_CFG2_SZ 32

`define GTYP_QUAD__CH0_ADAPT_LCK_CFG3    32'h00000024
`define GTYP_QUAD__CH0_ADAPT_LCK_CFG3_SZ 32

`define GTYP_QUAD__CH0_ADAPT_LOP_CFG    32'h00000025
`define GTYP_QUAD__CH0_ADAPT_LOP_CFG_SZ 32

`define GTYP_QUAD__CH0_ADAPT_OS_CFG    32'h00000026
`define GTYP_QUAD__CH0_ADAPT_OS_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_ILO_CFG    32'h00000027
`define GTYP_QUAD__CH0_CHCLK_ILO_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_MISC_CFG    32'h00000028
`define GTYP_QUAD__CH0_CHCLK_MISC_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_RSV_CFG    32'h00000029
`define GTYP_QUAD__CH0_CHCLK_RSV_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG    32'h0000002a
`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG1    32'h0000002b
`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG1_SZ 32

`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG2    32'h0000002c
`define GTYP_QUAD__CH0_CHCLK_RXCAL_CFG2_SZ 32

`define GTYP_QUAD__CH0_CHCLK_RXPI_CFG    32'h0000002d
`define GTYP_QUAD__CH0_CHCLK_RXPI_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_TXCAL_CFG    32'h0000002e
`define GTYP_QUAD__CH0_CHCLK_TXCAL_CFG_SZ 32

`define GTYP_QUAD__CH0_CHCLK_TXPI_CFG0    32'h0000002f
`define GTYP_QUAD__CH0_CHCLK_TXPI_CFG0_SZ 32

`define GTYP_QUAD__CH0_CHL_RSV_CFG0    32'h00000030
`define GTYP_QUAD__CH0_CHL_RSV_CFG0_SZ 32

`define GTYP_QUAD__CH0_CHL_RSV_CFG1    32'h00000031
`define GTYP_QUAD__CH0_CHL_RSV_CFG1_SZ 32

`define GTYP_QUAD__CH0_CHL_RSV_CFG2    32'h00000032
`define GTYP_QUAD__CH0_CHL_RSV_CFG2_SZ 32

`define GTYP_QUAD__CH0_CHL_RSV_CFG3    32'h00000033
`define GTYP_QUAD__CH0_CHL_RSV_CFG3_SZ 32

`define GTYP_QUAD__CH0_CHL_RSV_CFG4    32'h00000034
`define GTYP_QUAD__CH0_CHL_RSV_CFG4_SZ 32

`define GTYP_QUAD__CH0_DA_CFG    32'h00000035
`define GTYP_QUAD__CH0_DA_CFG_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG0    32'h00000036
`define GTYP_QUAD__CH0_EYESCAN_CFG0_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG1    32'h00000037
`define GTYP_QUAD__CH0_EYESCAN_CFG1_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG10    32'h00000038
`define GTYP_QUAD__CH0_EYESCAN_CFG10_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG11    32'h00000039
`define GTYP_QUAD__CH0_EYESCAN_CFG11_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG12    32'h0000003a
`define GTYP_QUAD__CH0_EYESCAN_CFG12_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG13    32'h0000003b
`define GTYP_QUAD__CH0_EYESCAN_CFG13_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG14    32'h0000003c
`define GTYP_QUAD__CH0_EYESCAN_CFG14_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG15    32'h0000003d
`define GTYP_QUAD__CH0_EYESCAN_CFG15_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG16    32'h0000003e
`define GTYP_QUAD__CH0_EYESCAN_CFG16_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG2    32'h0000003f
`define GTYP_QUAD__CH0_EYESCAN_CFG2_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG3    32'h00000040
`define GTYP_QUAD__CH0_EYESCAN_CFG3_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG4    32'h00000041
`define GTYP_QUAD__CH0_EYESCAN_CFG4_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG5    32'h00000042
`define GTYP_QUAD__CH0_EYESCAN_CFG5_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG6    32'h00000043
`define GTYP_QUAD__CH0_EYESCAN_CFG6_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG7    32'h00000044
`define GTYP_QUAD__CH0_EYESCAN_CFG7_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG8    32'h00000045
`define GTYP_QUAD__CH0_EYESCAN_CFG8_SZ 32

`define GTYP_QUAD__CH0_EYESCAN_CFG9    32'h00000046
`define GTYP_QUAD__CH0_EYESCAN_CFG9_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG0    32'h00000047
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG0_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG1    32'h00000048
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG1_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG2    32'h00000049
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG2_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG3    32'h0000004a
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG3_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG4    32'h0000004b
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG4_SZ 32

`define GTYP_QUAD__CH0_FABRIC_INTF_CFG5    32'h0000004c
`define GTYP_QUAD__CH0_FABRIC_INTF_CFG5_SZ 32

`define GTYP_QUAD__CH0_INSTANTIATED    32'h0000004d
`define GTYP_QUAD__CH0_INSTANTIATED_SZ 1

`define GTYP_QUAD__CH0_MONITOR_CFG    32'h0000004e
`define GTYP_QUAD__CH0_MONITOR_CFG_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG0    32'h0000004f
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG0_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG1    32'h00000050
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG1_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG10    32'h00000051
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG10_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG2    32'h00000052
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG2_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG3    32'h00000053
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG3_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG4    32'h00000054
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG4_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG5    32'h00000055
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG5_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG6    32'h00000056
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG6_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG7    32'h00000057
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG7_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG8    32'h00000058
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG8_SZ 32

`define GTYP_QUAD__CH0_PIPE_CTRL_CFG9    32'h00000059
`define GTYP_QUAD__CH0_PIPE_CTRL_CFG9_SZ 32

`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG0    32'h0000005a
`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG0_SZ 32

`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG1    32'h0000005b
`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG1_SZ 32

`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG2    32'h0000005c
`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG2_SZ 32

`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG3    32'h0000005d
`define GTYP_QUAD__CH0_PIPE_TX_EQ_CFG3_SZ 32

`define GTYP_QUAD__CH0_RESET_BYP_HDSHK_CFG    32'h0000005e
`define GTYP_QUAD__CH0_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYP_QUAD__CH0_RESET_CFG    32'h0000005f
`define GTYP_QUAD__CH0_RESET_CFG_SZ 32

`define GTYP_QUAD__CH0_RESET_LOOPER_ID_CFG    32'h00000060
`define GTYP_QUAD__CH0_RESET_LOOPER_ID_CFG_SZ 32

`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG0    32'h00000061
`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG0_SZ 32

`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG1    32'h00000062
`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG1_SZ 32

`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG2    32'h00000063
`define GTYP_QUAD__CH0_RESET_LOOP_ID_CFG2_SZ 32

`define GTYP_QUAD__CH0_RESET_TIME_CFG0    32'h00000064
`define GTYP_QUAD__CH0_RESET_TIME_CFG0_SZ 32

`define GTYP_QUAD__CH0_RESET_TIME_CFG1    32'h00000065
`define GTYP_QUAD__CH0_RESET_TIME_CFG1_SZ 32

`define GTYP_QUAD__CH0_RESET_TIME_CFG2    32'h00000066
`define GTYP_QUAD__CH0_RESET_TIME_CFG2_SZ 32

`define GTYP_QUAD__CH0_RESET_TIME_CFG3    32'h00000067
`define GTYP_QUAD__CH0_RESET_TIME_CFG3_SZ 32

`define GTYP_QUAD__CH0_RXOUTCLK_FREQ    32'h00000068
`define GTYP_QUAD__CH0_RXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH0_RXOUTCLK_REF_FREQ    32'h00000069
`define GTYP_QUAD__CH0_RXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH0_RXOUTCLK_REF_SOURCE    32'h0000006a
`define GTYP_QUAD__CH0_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH0_RX_CDR_CFG0    32'h0000006b
`define GTYP_QUAD__CH0_RX_CDR_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_CDR_CFG1    32'h0000006c
`define GTYP_QUAD__CH0_RX_CDR_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_CDR_CFG2    32'h0000006d
`define GTYP_QUAD__CH0_RX_CDR_CFG2_SZ 32

`define GTYP_QUAD__CH0_RX_CDR_CFG3    32'h0000006e
`define GTYP_QUAD__CH0_RX_CDR_CFG3_SZ 32

`define GTYP_QUAD__CH0_RX_CDR_CFG4    32'h0000006f
`define GTYP_QUAD__CH0_RX_CDR_CFG4_SZ 32

`define GTYP_QUAD__CH0_RX_CRC_CFG0    32'h00000070
`define GTYP_QUAD__CH0_RX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_CRC_CFG1    32'h00000071
`define GTYP_QUAD__CH0_RX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_CRC_CFG2    32'h00000072
`define GTYP_QUAD__CH0_RX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH0_RX_CRC_CFG3    32'h00000073
`define GTYP_QUAD__CH0_RX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH0_RX_CTLE_CFG0    32'h00000074
`define GTYP_QUAD__CH0_RX_CTLE_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_CTLE_CFG1    32'h00000075
`define GTYP_QUAD__CH0_RX_CTLE_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_DACI2V_CFG0    32'h00000076
`define GTYP_QUAD__CH0_RX_DACI2V_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_DATA_RATE    32'h00000077
`define GTYP_QUAD__CH0_RX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH0_RX_DFE_CFG0    32'h00000078
`define GTYP_QUAD__CH0_RX_DFE_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG0    32'h00000079
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG1    32'h0000007a
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG2    32'h0000007b
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG3    32'h0000007c
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG4    32'h0000007d
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG5    32'h0000007e
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG6    32'h0000007f
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG7    32'h00000080
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG8    32'h00000081
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG9    32'h00000082
`define GTYP_QUAD__CH0_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYP_QUAD__CH0_RX_MISC_CFG0    32'h00000083
`define GTYP_QUAD__CH0_RX_MISC_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_OOB_CFG0    32'h00000084
`define GTYP_QUAD__CH0_RX_OOB_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_OOB_CFG1    32'h00000085
`define GTYP_QUAD__CH0_RX_OOB_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_PAD_CFG0    32'h00000086
`define GTYP_QUAD__CH0_RX_PAD_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_PAD_CFG1    32'h00000087
`define GTYP_QUAD__CH0_RX_PAD_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_PCS_CFG0    32'h00000088
`define GTYP_QUAD__CH0_RX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_PCS_CFG1    32'h00000089
`define GTYP_QUAD__CH0_RX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_PCS_CFG2    32'h0000008a
`define GTYP_QUAD__CH0_RX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH0_RX_PCS_CFG3    32'h0000008b
`define GTYP_QUAD__CH0_RX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH0_RX_PCS_CFG4    32'h0000008c
`define GTYP_QUAD__CH0_RX_PCS_CFG4_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG0    32'h0000008d
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG1    32'h0000008e
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG2    32'h0000008f
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG3    32'h00000090
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG4    32'h00000091
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH0_RX_PHALIGN_CFG5    32'h00000092
`define GTYP_QUAD__CH0_RX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH0_SIM_MODE    32'h00000093
`define GTYP_QUAD__CH0_SIM_MODE_SZ 48

`define GTYP_QUAD__CH0_SIM_RECEIVER_DETECT_PASS    32'h00000094
`define GTYP_QUAD__CH0_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYP_QUAD__CH0_SIM_RESET_SPEEDUP    32'h00000095
`define GTYP_QUAD__CH0_SIM_RESET_SPEEDUP_SZ 40

`define GTYP_QUAD__CH0_SIM_TX_EIDLE_DRIVE_LEVEL    32'h00000096
`define GTYP_QUAD__CH0_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYP_QUAD__CH0_TXOUTCLK_FREQ    32'h00000097
`define GTYP_QUAD__CH0_TXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH0_TXOUTCLK_REF_FREQ    32'h00000098
`define GTYP_QUAD__CH0_TXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH0_TXOUTCLK_REF_SOURCE    32'h00000099
`define GTYP_QUAD__CH0_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH0_TX_10G_CFG0    32'h0000009a
`define GTYP_QUAD__CH0_TX_10G_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_10G_CFG1    32'h0000009b
`define GTYP_QUAD__CH0_TX_10G_CFG1_SZ 32

`define GTYP_QUAD__CH0_TX_10G_CFG2    32'h0000009c
`define GTYP_QUAD__CH0_TX_10G_CFG2_SZ 32

`define GTYP_QUAD__CH0_TX_10G_CFG3    32'h0000009d
`define GTYP_QUAD__CH0_TX_10G_CFG3_SZ 32

`define GTYP_QUAD__CH0_TX_ANA_CFG0    32'h0000009e
`define GTYP_QUAD__CH0_TX_ANA_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_CRC_CFG0    32'h0000009f
`define GTYP_QUAD__CH0_TX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_CRC_CFG1    32'h000000a0
`define GTYP_QUAD__CH0_TX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH0_TX_CRC_CFG2    32'h000000a1
`define GTYP_QUAD__CH0_TX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH0_TX_CRC_CFG3    32'h000000a2
`define GTYP_QUAD__CH0_TX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH0_TX_DATA_RATE    32'h000000a3
`define GTYP_QUAD__CH0_TX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH0_TX_DRV_CFG0    32'h000000a4
`define GTYP_QUAD__CH0_TX_DRV_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_DRV_CFG1    32'h000000a5
`define GTYP_QUAD__CH0_TX_DRV_CFG1_SZ 32

`define GTYP_QUAD__CH0_TX_PCS_CFG0    32'h000000a6
`define GTYP_QUAD__CH0_TX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_PCS_CFG1    32'h000000a7
`define GTYP_QUAD__CH0_TX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH0_TX_PCS_CFG2    32'h000000a8
`define GTYP_QUAD__CH0_TX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH0_TX_PCS_CFG3    32'h000000a9
`define GTYP_QUAD__CH0_TX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG0    32'h000000aa
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG1    32'h000000ab
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG2    32'h000000ac
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG3    32'h000000ad
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG4    32'h000000ae
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH0_TX_PHALIGN_CFG5    32'h000000af
`define GTYP_QUAD__CH0_TX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH0_TX_PIPPM_CFG    32'h000000b0
`define GTYP_QUAD__CH0_TX_PIPPM_CFG_SZ 32

`define GTYP_QUAD__CH0_TX_SER_CFG0    32'h000000b1
`define GTYP_QUAD__CH0_TX_SER_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_APT_CFG    32'h000000b2
`define GTYP_QUAD__CH1_ADAPT_APT_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_CAL_CFG    32'h000000b3
`define GTYP_QUAD__CH1_ADAPT_CAL_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_DFE_CFG    32'h000000b4
`define GTYP_QUAD__CH1_ADAPT_DFE_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GC_CFG0    32'h000000b5
`define GTYP_QUAD__CH1_ADAPT_GC_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GC_CFG1    32'h000000b6
`define GTYP_QUAD__CH1_ADAPT_GC_CFG1_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GC_CFG2    32'h000000b7
`define GTYP_QUAD__CH1_ADAPT_GC_CFG2_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GC_CFG3    32'h000000b8
`define GTYP_QUAD__CH1_ADAPT_GC_CFG3_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GEN_CFG0    32'h000000b9
`define GTYP_QUAD__CH1_ADAPT_GEN_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GEN_CFG1    32'h000000ba
`define GTYP_QUAD__CH1_ADAPT_GEN_CFG1_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GEN_CFG2    32'h000000bb
`define GTYP_QUAD__CH1_ADAPT_GEN_CFG2_SZ 32

`define GTYP_QUAD__CH1_ADAPT_GEN_CFG3    32'h000000bc
`define GTYP_QUAD__CH1_ADAPT_GEN_CFG3_SZ 32

`define GTYP_QUAD__CH1_ADAPT_H01_CFG    32'h000000bd
`define GTYP_QUAD__CH1_ADAPT_H01_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_H23_CFG    32'h000000be
`define GTYP_QUAD__CH1_ADAPT_H23_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_H45_CFG    32'h000000bf
`define GTYP_QUAD__CH1_ADAPT_H45_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_H67_CFG    32'h000000c0
`define GTYP_QUAD__CH1_ADAPT_H67_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_H89_CFG    32'h000000c1
`define GTYP_QUAD__CH1_ADAPT_H89_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_HAB_CFG    32'h000000c2
`define GTYP_QUAD__CH1_ADAPT_HAB_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_HCD_CFG    32'h000000c3
`define GTYP_QUAD__CH1_ADAPT_HCD_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_HEF_CFG    32'h000000c4
`define GTYP_QUAD__CH1_ADAPT_HEF_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG0    32'h000000c5
`define GTYP_QUAD__CH1_ADAPT_KH_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG1    32'h000000c6
`define GTYP_QUAD__CH1_ADAPT_KH_CFG1_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG2    32'h000000c7
`define GTYP_QUAD__CH1_ADAPT_KH_CFG2_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG3    32'h000000c8
`define GTYP_QUAD__CH1_ADAPT_KH_CFG3_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG4    32'h000000c9
`define GTYP_QUAD__CH1_ADAPT_KH_CFG4_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KH_CFG5    32'h000000ca
`define GTYP_QUAD__CH1_ADAPT_KH_CFG5_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KL_CFG0    32'h000000cb
`define GTYP_QUAD__CH1_ADAPT_KL_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_KL_CFG1    32'h000000cc
`define GTYP_QUAD__CH1_ADAPT_KL_CFG1_SZ 32

`define GTYP_QUAD__CH1_ADAPT_LCK_CFG0    32'h000000cd
`define GTYP_QUAD__CH1_ADAPT_LCK_CFG0_SZ 32

`define GTYP_QUAD__CH1_ADAPT_LCK_CFG1    32'h000000ce
`define GTYP_QUAD__CH1_ADAPT_LCK_CFG1_SZ 32

`define GTYP_QUAD__CH1_ADAPT_LCK_CFG2    32'h000000cf
`define GTYP_QUAD__CH1_ADAPT_LCK_CFG2_SZ 32

`define GTYP_QUAD__CH1_ADAPT_LCK_CFG3    32'h000000d0
`define GTYP_QUAD__CH1_ADAPT_LCK_CFG3_SZ 32

`define GTYP_QUAD__CH1_ADAPT_LOP_CFG    32'h000000d1
`define GTYP_QUAD__CH1_ADAPT_LOP_CFG_SZ 32

`define GTYP_QUAD__CH1_ADAPT_OS_CFG    32'h000000d2
`define GTYP_QUAD__CH1_ADAPT_OS_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_ILO_CFG    32'h000000d3
`define GTYP_QUAD__CH1_CHCLK_ILO_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_MISC_CFG    32'h000000d4
`define GTYP_QUAD__CH1_CHCLK_MISC_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_RSV_CFG    32'h000000d5
`define GTYP_QUAD__CH1_CHCLK_RSV_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG    32'h000000d6
`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG1    32'h000000d7
`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG1_SZ 32

`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG2    32'h000000d8
`define GTYP_QUAD__CH1_CHCLK_RXCAL_CFG2_SZ 32

`define GTYP_QUAD__CH1_CHCLK_RXPI_CFG    32'h000000d9
`define GTYP_QUAD__CH1_CHCLK_RXPI_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_TXCAL_CFG    32'h000000da
`define GTYP_QUAD__CH1_CHCLK_TXCAL_CFG_SZ 32

`define GTYP_QUAD__CH1_CHCLK_TXPI_CFG0    32'h000000db
`define GTYP_QUAD__CH1_CHCLK_TXPI_CFG0_SZ 32

`define GTYP_QUAD__CH1_CHL_RSV_CFG0    32'h000000dc
`define GTYP_QUAD__CH1_CHL_RSV_CFG0_SZ 32

`define GTYP_QUAD__CH1_CHL_RSV_CFG1    32'h000000dd
`define GTYP_QUAD__CH1_CHL_RSV_CFG1_SZ 32

`define GTYP_QUAD__CH1_CHL_RSV_CFG2    32'h000000de
`define GTYP_QUAD__CH1_CHL_RSV_CFG2_SZ 32

`define GTYP_QUAD__CH1_CHL_RSV_CFG3    32'h000000df
`define GTYP_QUAD__CH1_CHL_RSV_CFG3_SZ 32

`define GTYP_QUAD__CH1_CHL_RSV_CFG4    32'h000000e0
`define GTYP_QUAD__CH1_CHL_RSV_CFG4_SZ 32

`define GTYP_QUAD__CH1_DA_CFG    32'h000000e1
`define GTYP_QUAD__CH1_DA_CFG_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG0    32'h000000e2
`define GTYP_QUAD__CH1_EYESCAN_CFG0_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG1    32'h000000e3
`define GTYP_QUAD__CH1_EYESCAN_CFG1_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG10    32'h000000e4
`define GTYP_QUAD__CH1_EYESCAN_CFG10_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG11    32'h000000e5
`define GTYP_QUAD__CH1_EYESCAN_CFG11_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG12    32'h000000e6
`define GTYP_QUAD__CH1_EYESCAN_CFG12_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG13    32'h000000e7
`define GTYP_QUAD__CH1_EYESCAN_CFG13_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG14    32'h000000e8
`define GTYP_QUAD__CH1_EYESCAN_CFG14_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG15    32'h000000e9
`define GTYP_QUAD__CH1_EYESCAN_CFG15_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG16    32'h000000ea
`define GTYP_QUAD__CH1_EYESCAN_CFG16_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG2    32'h000000eb
`define GTYP_QUAD__CH1_EYESCAN_CFG2_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG3    32'h000000ec
`define GTYP_QUAD__CH1_EYESCAN_CFG3_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG4    32'h000000ed
`define GTYP_QUAD__CH1_EYESCAN_CFG4_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG5    32'h000000ee
`define GTYP_QUAD__CH1_EYESCAN_CFG5_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG6    32'h000000ef
`define GTYP_QUAD__CH1_EYESCAN_CFG6_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG7    32'h000000f0
`define GTYP_QUAD__CH1_EYESCAN_CFG7_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG8    32'h000000f1
`define GTYP_QUAD__CH1_EYESCAN_CFG8_SZ 32

`define GTYP_QUAD__CH1_EYESCAN_CFG9    32'h000000f2
`define GTYP_QUAD__CH1_EYESCAN_CFG9_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG0    32'h000000f3
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG0_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG1    32'h000000f4
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG1_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG2    32'h000000f5
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG2_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG3    32'h000000f6
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG3_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG4    32'h000000f7
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG4_SZ 32

`define GTYP_QUAD__CH1_FABRIC_INTF_CFG5    32'h000000f8
`define GTYP_QUAD__CH1_FABRIC_INTF_CFG5_SZ 32

`define GTYP_QUAD__CH1_INSTANTIATED    32'h000000f9
`define GTYP_QUAD__CH1_INSTANTIATED_SZ 1

`define GTYP_QUAD__CH1_MONITOR_CFG    32'h000000fa
`define GTYP_QUAD__CH1_MONITOR_CFG_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG0    32'h000000fb
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG0_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG1    32'h000000fc
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG1_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG10    32'h000000fd
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG10_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG2    32'h000000fe
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG2_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG3    32'h000000ff
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG3_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG4    32'h00000100
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG4_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG5    32'h00000101
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG5_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG6    32'h00000102
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG6_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG7    32'h00000103
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG7_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG8    32'h00000104
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG8_SZ 32

`define GTYP_QUAD__CH1_PIPE_CTRL_CFG9    32'h00000105
`define GTYP_QUAD__CH1_PIPE_CTRL_CFG9_SZ 32

`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG0    32'h00000106
`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG0_SZ 32

`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG1    32'h00000107
`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG1_SZ 32

`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG2    32'h00000108
`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG2_SZ 32

`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG3    32'h00000109
`define GTYP_QUAD__CH1_PIPE_TX_EQ_CFG3_SZ 32

`define GTYP_QUAD__CH1_RESET_BYP_HDSHK_CFG    32'h0000010a
`define GTYP_QUAD__CH1_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYP_QUAD__CH1_RESET_CFG    32'h0000010b
`define GTYP_QUAD__CH1_RESET_CFG_SZ 32

`define GTYP_QUAD__CH1_RESET_LOOPER_ID_CFG    32'h0000010c
`define GTYP_QUAD__CH1_RESET_LOOPER_ID_CFG_SZ 32

`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG0    32'h0000010d
`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG0_SZ 32

`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG1    32'h0000010e
`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG1_SZ 32

`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG2    32'h0000010f
`define GTYP_QUAD__CH1_RESET_LOOP_ID_CFG2_SZ 32

`define GTYP_QUAD__CH1_RESET_TIME_CFG0    32'h00000110
`define GTYP_QUAD__CH1_RESET_TIME_CFG0_SZ 32

`define GTYP_QUAD__CH1_RESET_TIME_CFG1    32'h00000111
`define GTYP_QUAD__CH1_RESET_TIME_CFG1_SZ 32

`define GTYP_QUAD__CH1_RESET_TIME_CFG2    32'h00000112
`define GTYP_QUAD__CH1_RESET_TIME_CFG2_SZ 32

`define GTYP_QUAD__CH1_RESET_TIME_CFG3    32'h00000113
`define GTYP_QUAD__CH1_RESET_TIME_CFG3_SZ 32

`define GTYP_QUAD__CH1_RXOUTCLK_FREQ    32'h00000114
`define GTYP_QUAD__CH1_RXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH1_RXOUTCLK_REF_FREQ    32'h00000115
`define GTYP_QUAD__CH1_RXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH1_RXOUTCLK_REF_SOURCE    32'h00000116
`define GTYP_QUAD__CH1_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH1_RX_CDR_CFG0    32'h00000117
`define GTYP_QUAD__CH1_RX_CDR_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_CDR_CFG1    32'h00000118
`define GTYP_QUAD__CH1_RX_CDR_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_CDR_CFG2    32'h00000119
`define GTYP_QUAD__CH1_RX_CDR_CFG2_SZ 32

`define GTYP_QUAD__CH1_RX_CDR_CFG3    32'h0000011a
`define GTYP_QUAD__CH1_RX_CDR_CFG3_SZ 32

`define GTYP_QUAD__CH1_RX_CDR_CFG4    32'h0000011b
`define GTYP_QUAD__CH1_RX_CDR_CFG4_SZ 32

`define GTYP_QUAD__CH1_RX_CRC_CFG0    32'h0000011c
`define GTYP_QUAD__CH1_RX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_CRC_CFG1    32'h0000011d
`define GTYP_QUAD__CH1_RX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_CRC_CFG2    32'h0000011e
`define GTYP_QUAD__CH1_RX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH1_RX_CRC_CFG3    32'h0000011f
`define GTYP_QUAD__CH1_RX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH1_RX_CTLE_CFG0    32'h00000120
`define GTYP_QUAD__CH1_RX_CTLE_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_CTLE_CFG1    32'h00000121
`define GTYP_QUAD__CH1_RX_CTLE_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_DACI2V_CFG0    32'h00000122
`define GTYP_QUAD__CH1_RX_DACI2V_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_DATA_RATE    32'h00000123
`define GTYP_QUAD__CH1_RX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH1_RX_DFE_CFG0    32'h00000124
`define GTYP_QUAD__CH1_RX_DFE_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG0    32'h00000125
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG1    32'h00000126
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG2    32'h00000127
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG3    32'h00000128
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG4    32'h00000129
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG5    32'h0000012a
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG6    32'h0000012b
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG7    32'h0000012c
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG8    32'h0000012d
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG9    32'h0000012e
`define GTYP_QUAD__CH1_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYP_QUAD__CH1_RX_MISC_CFG0    32'h0000012f
`define GTYP_QUAD__CH1_RX_MISC_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_OOB_CFG0    32'h00000130
`define GTYP_QUAD__CH1_RX_OOB_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_OOB_CFG1    32'h00000131
`define GTYP_QUAD__CH1_RX_OOB_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_PAD_CFG0    32'h00000132
`define GTYP_QUAD__CH1_RX_PAD_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_PAD_CFG1    32'h00000133
`define GTYP_QUAD__CH1_RX_PAD_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_PCS_CFG0    32'h00000134
`define GTYP_QUAD__CH1_RX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_PCS_CFG1    32'h00000135
`define GTYP_QUAD__CH1_RX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_PCS_CFG2    32'h00000136
`define GTYP_QUAD__CH1_RX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH1_RX_PCS_CFG3    32'h00000137
`define GTYP_QUAD__CH1_RX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH1_RX_PCS_CFG4    32'h00000138
`define GTYP_QUAD__CH1_RX_PCS_CFG4_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG0    32'h00000139
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG1    32'h0000013a
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG2    32'h0000013b
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG3    32'h0000013c
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG4    32'h0000013d
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH1_RX_PHALIGN_CFG5    32'h0000013e
`define GTYP_QUAD__CH1_RX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH1_SIM_MODE    32'h0000013f
`define GTYP_QUAD__CH1_SIM_MODE_SZ 48

`define GTYP_QUAD__CH1_SIM_RECEIVER_DETECT_PASS    32'h00000140
`define GTYP_QUAD__CH1_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYP_QUAD__CH1_SIM_RESET_SPEEDUP    32'h00000141
`define GTYP_QUAD__CH1_SIM_RESET_SPEEDUP_SZ 40

`define GTYP_QUAD__CH1_SIM_TX_EIDLE_DRIVE_LEVEL    32'h00000142
`define GTYP_QUAD__CH1_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYP_QUAD__CH1_TXOUTCLK_FREQ    32'h00000143
`define GTYP_QUAD__CH1_TXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH1_TXOUTCLK_REF_FREQ    32'h00000144
`define GTYP_QUAD__CH1_TXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH1_TXOUTCLK_REF_SOURCE    32'h00000145
`define GTYP_QUAD__CH1_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH1_TX_10G_CFG0    32'h00000146
`define GTYP_QUAD__CH1_TX_10G_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_10G_CFG1    32'h00000147
`define GTYP_QUAD__CH1_TX_10G_CFG1_SZ 32

`define GTYP_QUAD__CH1_TX_10G_CFG2    32'h00000148
`define GTYP_QUAD__CH1_TX_10G_CFG2_SZ 32

`define GTYP_QUAD__CH1_TX_10G_CFG3    32'h00000149
`define GTYP_QUAD__CH1_TX_10G_CFG3_SZ 32

`define GTYP_QUAD__CH1_TX_ANA_CFG0    32'h0000014a
`define GTYP_QUAD__CH1_TX_ANA_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_CRC_CFG0    32'h0000014b
`define GTYP_QUAD__CH1_TX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_CRC_CFG1    32'h0000014c
`define GTYP_QUAD__CH1_TX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH1_TX_CRC_CFG2    32'h0000014d
`define GTYP_QUAD__CH1_TX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH1_TX_CRC_CFG3    32'h0000014e
`define GTYP_QUAD__CH1_TX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH1_TX_DATA_RATE    32'h0000014f
`define GTYP_QUAD__CH1_TX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH1_TX_DRV_CFG0    32'h00000150
`define GTYP_QUAD__CH1_TX_DRV_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_DRV_CFG1    32'h00000151
`define GTYP_QUAD__CH1_TX_DRV_CFG1_SZ 32

`define GTYP_QUAD__CH1_TX_PCS_CFG0    32'h00000152
`define GTYP_QUAD__CH1_TX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_PCS_CFG1    32'h00000153
`define GTYP_QUAD__CH1_TX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH1_TX_PCS_CFG2    32'h00000154
`define GTYP_QUAD__CH1_TX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH1_TX_PCS_CFG3    32'h00000155
`define GTYP_QUAD__CH1_TX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG0    32'h00000156
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG1    32'h00000157
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG2    32'h00000158
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG3    32'h00000159
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG4    32'h0000015a
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH1_TX_PHALIGN_CFG5    32'h0000015b
`define GTYP_QUAD__CH1_TX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH1_TX_PIPPM_CFG    32'h0000015c
`define GTYP_QUAD__CH1_TX_PIPPM_CFG_SZ 32

`define GTYP_QUAD__CH1_TX_SER_CFG0    32'h0000015d
`define GTYP_QUAD__CH1_TX_SER_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_APT_CFG    32'h0000015e
`define GTYP_QUAD__CH2_ADAPT_APT_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_CAL_CFG    32'h0000015f
`define GTYP_QUAD__CH2_ADAPT_CAL_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_DFE_CFG    32'h00000160
`define GTYP_QUAD__CH2_ADAPT_DFE_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GC_CFG0    32'h00000161
`define GTYP_QUAD__CH2_ADAPT_GC_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GC_CFG1    32'h00000162
`define GTYP_QUAD__CH2_ADAPT_GC_CFG1_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GC_CFG2    32'h00000163
`define GTYP_QUAD__CH2_ADAPT_GC_CFG2_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GC_CFG3    32'h00000164
`define GTYP_QUAD__CH2_ADAPT_GC_CFG3_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GEN_CFG0    32'h00000165
`define GTYP_QUAD__CH2_ADAPT_GEN_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GEN_CFG1    32'h00000166
`define GTYP_QUAD__CH2_ADAPT_GEN_CFG1_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GEN_CFG2    32'h00000167
`define GTYP_QUAD__CH2_ADAPT_GEN_CFG2_SZ 32

`define GTYP_QUAD__CH2_ADAPT_GEN_CFG3    32'h00000168
`define GTYP_QUAD__CH2_ADAPT_GEN_CFG3_SZ 32

`define GTYP_QUAD__CH2_ADAPT_H01_CFG    32'h00000169
`define GTYP_QUAD__CH2_ADAPT_H01_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_H23_CFG    32'h0000016a
`define GTYP_QUAD__CH2_ADAPT_H23_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_H45_CFG    32'h0000016b
`define GTYP_QUAD__CH2_ADAPT_H45_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_H67_CFG    32'h0000016c
`define GTYP_QUAD__CH2_ADAPT_H67_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_H89_CFG    32'h0000016d
`define GTYP_QUAD__CH2_ADAPT_H89_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_HAB_CFG    32'h0000016e
`define GTYP_QUAD__CH2_ADAPT_HAB_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_HCD_CFG    32'h0000016f
`define GTYP_QUAD__CH2_ADAPT_HCD_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_HEF_CFG    32'h00000170
`define GTYP_QUAD__CH2_ADAPT_HEF_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG0    32'h00000171
`define GTYP_QUAD__CH2_ADAPT_KH_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG1    32'h00000172
`define GTYP_QUAD__CH2_ADAPT_KH_CFG1_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG2    32'h00000173
`define GTYP_QUAD__CH2_ADAPT_KH_CFG2_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG3    32'h00000174
`define GTYP_QUAD__CH2_ADAPT_KH_CFG3_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG4    32'h00000175
`define GTYP_QUAD__CH2_ADAPT_KH_CFG4_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KH_CFG5    32'h00000176
`define GTYP_QUAD__CH2_ADAPT_KH_CFG5_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KL_CFG0    32'h00000177
`define GTYP_QUAD__CH2_ADAPT_KL_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_KL_CFG1    32'h00000178
`define GTYP_QUAD__CH2_ADAPT_KL_CFG1_SZ 32

`define GTYP_QUAD__CH2_ADAPT_LCK_CFG0    32'h00000179
`define GTYP_QUAD__CH2_ADAPT_LCK_CFG0_SZ 32

`define GTYP_QUAD__CH2_ADAPT_LCK_CFG1    32'h0000017a
`define GTYP_QUAD__CH2_ADAPT_LCK_CFG1_SZ 32

`define GTYP_QUAD__CH2_ADAPT_LCK_CFG2    32'h0000017b
`define GTYP_QUAD__CH2_ADAPT_LCK_CFG2_SZ 32

`define GTYP_QUAD__CH2_ADAPT_LCK_CFG3    32'h0000017c
`define GTYP_QUAD__CH2_ADAPT_LCK_CFG3_SZ 32

`define GTYP_QUAD__CH2_ADAPT_LOP_CFG    32'h0000017d
`define GTYP_QUAD__CH2_ADAPT_LOP_CFG_SZ 32

`define GTYP_QUAD__CH2_ADAPT_OS_CFG    32'h0000017e
`define GTYP_QUAD__CH2_ADAPT_OS_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_ILO_CFG    32'h0000017f
`define GTYP_QUAD__CH2_CHCLK_ILO_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_MISC_CFG    32'h00000180
`define GTYP_QUAD__CH2_CHCLK_MISC_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_RSV_CFG    32'h00000181
`define GTYP_QUAD__CH2_CHCLK_RSV_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG    32'h00000182
`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG1    32'h00000183
`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG1_SZ 32

`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG2    32'h00000184
`define GTYP_QUAD__CH2_CHCLK_RXCAL_CFG2_SZ 32

`define GTYP_QUAD__CH2_CHCLK_RXPI_CFG    32'h00000185
`define GTYP_QUAD__CH2_CHCLK_RXPI_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_TXCAL_CFG    32'h00000186
`define GTYP_QUAD__CH2_CHCLK_TXCAL_CFG_SZ 32

`define GTYP_QUAD__CH2_CHCLK_TXPI_CFG0    32'h00000187
`define GTYP_QUAD__CH2_CHCLK_TXPI_CFG0_SZ 32

`define GTYP_QUAD__CH2_CHL_RSV_CFG0    32'h00000188
`define GTYP_QUAD__CH2_CHL_RSV_CFG0_SZ 32

`define GTYP_QUAD__CH2_CHL_RSV_CFG1    32'h00000189
`define GTYP_QUAD__CH2_CHL_RSV_CFG1_SZ 32

`define GTYP_QUAD__CH2_CHL_RSV_CFG2    32'h0000018a
`define GTYP_QUAD__CH2_CHL_RSV_CFG2_SZ 32

`define GTYP_QUAD__CH2_CHL_RSV_CFG3    32'h0000018b
`define GTYP_QUAD__CH2_CHL_RSV_CFG3_SZ 32

`define GTYP_QUAD__CH2_CHL_RSV_CFG4    32'h0000018c
`define GTYP_QUAD__CH2_CHL_RSV_CFG4_SZ 32

`define GTYP_QUAD__CH2_DA_CFG    32'h0000018d
`define GTYP_QUAD__CH2_DA_CFG_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG0    32'h0000018e
`define GTYP_QUAD__CH2_EYESCAN_CFG0_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG1    32'h0000018f
`define GTYP_QUAD__CH2_EYESCAN_CFG1_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG10    32'h00000190
`define GTYP_QUAD__CH2_EYESCAN_CFG10_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG11    32'h00000191
`define GTYP_QUAD__CH2_EYESCAN_CFG11_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG12    32'h00000192
`define GTYP_QUAD__CH2_EYESCAN_CFG12_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG13    32'h00000193
`define GTYP_QUAD__CH2_EYESCAN_CFG13_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG14    32'h00000194
`define GTYP_QUAD__CH2_EYESCAN_CFG14_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG15    32'h00000195
`define GTYP_QUAD__CH2_EYESCAN_CFG15_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG16    32'h00000196
`define GTYP_QUAD__CH2_EYESCAN_CFG16_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG2    32'h00000197
`define GTYP_QUAD__CH2_EYESCAN_CFG2_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG3    32'h00000198
`define GTYP_QUAD__CH2_EYESCAN_CFG3_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG4    32'h00000199
`define GTYP_QUAD__CH2_EYESCAN_CFG4_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG5    32'h0000019a
`define GTYP_QUAD__CH2_EYESCAN_CFG5_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG6    32'h0000019b
`define GTYP_QUAD__CH2_EYESCAN_CFG6_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG7    32'h0000019c
`define GTYP_QUAD__CH2_EYESCAN_CFG7_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG8    32'h0000019d
`define GTYP_QUAD__CH2_EYESCAN_CFG8_SZ 32

`define GTYP_QUAD__CH2_EYESCAN_CFG9    32'h0000019e
`define GTYP_QUAD__CH2_EYESCAN_CFG9_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG0    32'h0000019f
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG0_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG1    32'h000001a0
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG1_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG2    32'h000001a1
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG2_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG3    32'h000001a2
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG3_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG4    32'h000001a3
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG4_SZ 32

`define GTYP_QUAD__CH2_FABRIC_INTF_CFG5    32'h000001a4
`define GTYP_QUAD__CH2_FABRIC_INTF_CFG5_SZ 32

`define GTYP_QUAD__CH2_INSTANTIATED    32'h000001a5
`define GTYP_QUAD__CH2_INSTANTIATED_SZ 1

`define GTYP_QUAD__CH2_MONITOR_CFG    32'h000001a6
`define GTYP_QUAD__CH2_MONITOR_CFG_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG0    32'h000001a7
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG0_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG1    32'h000001a8
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG1_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG10    32'h000001a9
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG10_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG2    32'h000001aa
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG2_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG3    32'h000001ab
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG3_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG4    32'h000001ac
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG4_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG5    32'h000001ad
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG5_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG6    32'h000001ae
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG6_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG7    32'h000001af
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG7_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG8    32'h000001b0
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG8_SZ 32

`define GTYP_QUAD__CH2_PIPE_CTRL_CFG9    32'h000001b1
`define GTYP_QUAD__CH2_PIPE_CTRL_CFG9_SZ 32

`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG0    32'h000001b2
`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG0_SZ 32

`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG1    32'h000001b3
`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG1_SZ 32

`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG2    32'h000001b4
`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG2_SZ 32

`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG3    32'h000001b5
`define GTYP_QUAD__CH2_PIPE_TX_EQ_CFG3_SZ 32

`define GTYP_QUAD__CH2_RESET_BYP_HDSHK_CFG    32'h000001b6
`define GTYP_QUAD__CH2_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYP_QUAD__CH2_RESET_CFG    32'h000001b7
`define GTYP_QUAD__CH2_RESET_CFG_SZ 32

`define GTYP_QUAD__CH2_RESET_LOOPER_ID_CFG    32'h000001b8
`define GTYP_QUAD__CH2_RESET_LOOPER_ID_CFG_SZ 32

`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG0    32'h000001b9
`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG0_SZ 32

`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG1    32'h000001ba
`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG1_SZ 32

`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG2    32'h000001bb
`define GTYP_QUAD__CH2_RESET_LOOP_ID_CFG2_SZ 32

`define GTYP_QUAD__CH2_RESET_TIME_CFG0    32'h000001bc
`define GTYP_QUAD__CH2_RESET_TIME_CFG0_SZ 32

`define GTYP_QUAD__CH2_RESET_TIME_CFG1    32'h000001bd
`define GTYP_QUAD__CH2_RESET_TIME_CFG1_SZ 32

`define GTYP_QUAD__CH2_RESET_TIME_CFG2    32'h000001be
`define GTYP_QUAD__CH2_RESET_TIME_CFG2_SZ 32

`define GTYP_QUAD__CH2_RESET_TIME_CFG3    32'h000001bf
`define GTYP_QUAD__CH2_RESET_TIME_CFG3_SZ 32

`define GTYP_QUAD__CH2_RXOUTCLK_FREQ    32'h000001c0
`define GTYP_QUAD__CH2_RXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH2_RXOUTCLK_REF_FREQ    32'h000001c1
`define GTYP_QUAD__CH2_RXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH2_RXOUTCLK_REF_SOURCE    32'h000001c2
`define GTYP_QUAD__CH2_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH2_RX_CDR_CFG0    32'h000001c3
`define GTYP_QUAD__CH2_RX_CDR_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_CDR_CFG1    32'h000001c4
`define GTYP_QUAD__CH2_RX_CDR_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_CDR_CFG2    32'h000001c5
`define GTYP_QUAD__CH2_RX_CDR_CFG2_SZ 32

`define GTYP_QUAD__CH2_RX_CDR_CFG3    32'h000001c6
`define GTYP_QUAD__CH2_RX_CDR_CFG3_SZ 32

`define GTYP_QUAD__CH2_RX_CDR_CFG4    32'h000001c7
`define GTYP_QUAD__CH2_RX_CDR_CFG4_SZ 32

`define GTYP_QUAD__CH2_RX_CRC_CFG0    32'h000001c8
`define GTYP_QUAD__CH2_RX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_CRC_CFG1    32'h000001c9
`define GTYP_QUAD__CH2_RX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_CRC_CFG2    32'h000001ca
`define GTYP_QUAD__CH2_RX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH2_RX_CRC_CFG3    32'h000001cb
`define GTYP_QUAD__CH2_RX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH2_RX_CTLE_CFG0    32'h000001cc
`define GTYP_QUAD__CH2_RX_CTLE_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_CTLE_CFG1    32'h000001cd
`define GTYP_QUAD__CH2_RX_CTLE_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_DACI2V_CFG0    32'h000001ce
`define GTYP_QUAD__CH2_RX_DACI2V_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_DATA_RATE    32'h000001cf
`define GTYP_QUAD__CH2_RX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH2_RX_DFE_CFG0    32'h000001d0
`define GTYP_QUAD__CH2_RX_DFE_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG0    32'h000001d1
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG1    32'h000001d2
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG2    32'h000001d3
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG3    32'h000001d4
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG4    32'h000001d5
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG5    32'h000001d6
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG6    32'h000001d7
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG7    32'h000001d8
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG8    32'h000001d9
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG9    32'h000001da
`define GTYP_QUAD__CH2_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYP_QUAD__CH2_RX_MISC_CFG0    32'h000001db
`define GTYP_QUAD__CH2_RX_MISC_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_OOB_CFG0    32'h000001dc
`define GTYP_QUAD__CH2_RX_OOB_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_OOB_CFG1    32'h000001dd
`define GTYP_QUAD__CH2_RX_OOB_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_PAD_CFG0    32'h000001de
`define GTYP_QUAD__CH2_RX_PAD_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_PAD_CFG1    32'h000001df
`define GTYP_QUAD__CH2_RX_PAD_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_PCS_CFG0    32'h000001e0
`define GTYP_QUAD__CH2_RX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_PCS_CFG1    32'h000001e1
`define GTYP_QUAD__CH2_RX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_PCS_CFG2    32'h000001e2
`define GTYP_QUAD__CH2_RX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH2_RX_PCS_CFG3    32'h000001e3
`define GTYP_QUAD__CH2_RX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH2_RX_PCS_CFG4    32'h000001e4
`define GTYP_QUAD__CH2_RX_PCS_CFG4_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG0    32'h000001e5
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG1    32'h000001e6
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG2    32'h000001e7
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG3    32'h000001e8
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG4    32'h000001e9
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH2_RX_PHALIGN_CFG5    32'h000001ea
`define GTYP_QUAD__CH2_RX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH2_SIM_MODE    32'h000001eb
`define GTYP_QUAD__CH2_SIM_MODE_SZ 48

`define GTYP_QUAD__CH2_SIM_RECEIVER_DETECT_PASS    32'h000001ec
`define GTYP_QUAD__CH2_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYP_QUAD__CH2_SIM_RESET_SPEEDUP    32'h000001ed
`define GTYP_QUAD__CH2_SIM_RESET_SPEEDUP_SZ 40

`define GTYP_QUAD__CH2_SIM_TX_EIDLE_DRIVE_LEVEL    32'h000001ee
`define GTYP_QUAD__CH2_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYP_QUAD__CH2_TXOUTCLK_FREQ    32'h000001ef
`define GTYP_QUAD__CH2_TXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH2_TXOUTCLK_REF_FREQ    32'h000001f0
`define GTYP_QUAD__CH2_TXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH2_TXOUTCLK_REF_SOURCE    32'h000001f1
`define GTYP_QUAD__CH2_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH2_TX_10G_CFG0    32'h000001f2
`define GTYP_QUAD__CH2_TX_10G_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_10G_CFG1    32'h000001f3
`define GTYP_QUAD__CH2_TX_10G_CFG1_SZ 32

`define GTYP_QUAD__CH2_TX_10G_CFG2    32'h000001f4
`define GTYP_QUAD__CH2_TX_10G_CFG2_SZ 32

`define GTYP_QUAD__CH2_TX_10G_CFG3    32'h000001f5
`define GTYP_QUAD__CH2_TX_10G_CFG3_SZ 32

`define GTYP_QUAD__CH2_TX_ANA_CFG0    32'h000001f6
`define GTYP_QUAD__CH2_TX_ANA_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_CRC_CFG0    32'h000001f7
`define GTYP_QUAD__CH2_TX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_CRC_CFG1    32'h000001f8
`define GTYP_QUAD__CH2_TX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH2_TX_CRC_CFG2    32'h000001f9
`define GTYP_QUAD__CH2_TX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH2_TX_CRC_CFG3    32'h000001fa
`define GTYP_QUAD__CH2_TX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH2_TX_DATA_RATE    32'h000001fb
`define GTYP_QUAD__CH2_TX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH2_TX_DRV_CFG0    32'h000001fc
`define GTYP_QUAD__CH2_TX_DRV_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_DRV_CFG1    32'h000001fd
`define GTYP_QUAD__CH2_TX_DRV_CFG1_SZ 32

`define GTYP_QUAD__CH2_TX_PCS_CFG0    32'h000001fe
`define GTYP_QUAD__CH2_TX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_PCS_CFG1    32'h000001ff
`define GTYP_QUAD__CH2_TX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH2_TX_PCS_CFG2    32'h00000200
`define GTYP_QUAD__CH2_TX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH2_TX_PCS_CFG3    32'h00000201
`define GTYP_QUAD__CH2_TX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG0    32'h00000202
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG1    32'h00000203
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG2    32'h00000204
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG3    32'h00000205
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG4    32'h00000206
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH2_TX_PHALIGN_CFG5    32'h00000207
`define GTYP_QUAD__CH2_TX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH2_TX_PIPPM_CFG    32'h00000208
`define GTYP_QUAD__CH2_TX_PIPPM_CFG_SZ 32

`define GTYP_QUAD__CH2_TX_SER_CFG0    32'h00000209
`define GTYP_QUAD__CH2_TX_SER_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_APT_CFG    32'h0000020a
`define GTYP_QUAD__CH3_ADAPT_APT_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_CAL_CFG    32'h0000020b
`define GTYP_QUAD__CH3_ADAPT_CAL_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_DFE_CFG    32'h0000020c
`define GTYP_QUAD__CH3_ADAPT_DFE_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GC_CFG0    32'h0000020d
`define GTYP_QUAD__CH3_ADAPT_GC_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GC_CFG1    32'h0000020e
`define GTYP_QUAD__CH3_ADAPT_GC_CFG1_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GC_CFG2    32'h0000020f
`define GTYP_QUAD__CH3_ADAPT_GC_CFG2_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GC_CFG3    32'h00000210
`define GTYP_QUAD__CH3_ADAPT_GC_CFG3_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GEN_CFG0    32'h00000211
`define GTYP_QUAD__CH3_ADAPT_GEN_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GEN_CFG1    32'h00000212
`define GTYP_QUAD__CH3_ADAPT_GEN_CFG1_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GEN_CFG2    32'h00000213
`define GTYP_QUAD__CH3_ADAPT_GEN_CFG2_SZ 32

`define GTYP_QUAD__CH3_ADAPT_GEN_CFG3    32'h00000214
`define GTYP_QUAD__CH3_ADAPT_GEN_CFG3_SZ 32

`define GTYP_QUAD__CH3_ADAPT_H01_CFG    32'h00000215
`define GTYP_QUAD__CH3_ADAPT_H01_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_H23_CFG    32'h00000216
`define GTYP_QUAD__CH3_ADAPT_H23_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_H45_CFG    32'h00000217
`define GTYP_QUAD__CH3_ADAPT_H45_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_H67_CFG    32'h00000218
`define GTYP_QUAD__CH3_ADAPT_H67_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_H89_CFG    32'h00000219
`define GTYP_QUAD__CH3_ADAPT_H89_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_HAB_CFG    32'h0000021a
`define GTYP_QUAD__CH3_ADAPT_HAB_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_HCD_CFG    32'h0000021b
`define GTYP_QUAD__CH3_ADAPT_HCD_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_HEF_CFG    32'h0000021c
`define GTYP_QUAD__CH3_ADAPT_HEF_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG0    32'h0000021d
`define GTYP_QUAD__CH3_ADAPT_KH_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG1    32'h0000021e
`define GTYP_QUAD__CH3_ADAPT_KH_CFG1_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG2    32'h0000021f
`define GTYP_QUAD__CH3_ADAPT_KH_CFG2_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG3    32'h00000220
`define GTYP_QUAD__CH3_ADAPT_KH_CFG3_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG4    32'h00000221
`define GTYP_QUAD__CH3_ADAPT_KH_CFG4_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KH_CFG5    32'h00000222
`define GTYP_QUAD__CH3_ADAPT_KH_CFG5_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KL_CFG0    32'h00000223
`define GTYP_QUAD__CH3_ADAPT_KL_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_KL_CFG1    32'h00000224
`define GTYP_QUAD__CH3_ADAPT_KL_CFG1_SZ 32

`define GTYP_QUAD__CH3_ADAPT_LCK_CFG0    32'h00000225
`define GTYP_QUAD__CH3_ADAPT_LCK_CFG0_SZ 32

`define GTYP_QUAD__CH3_ADAPT_LCK_CFG1    32'h00000226
`define GTYP_QUAD__CH3_ADAPT_LCK_CFG1_SZ 32

`define GTYP_QUAD__CH3_ADAPT_LCK_CFG2    32'h00000227
`define GTYP_QUAD__CH3_ADAPT_LCK_CFG2_SZ 32

`define GTYP_QUAD__CH3_ADAPT_LCK_CFG3    32'h00000228
`define GTYP_QUAD__CH3_ADAPT_LCK_CFG3_SZ 32

`define GTYP_QUAD__CH3_ADAPT_LOP_CFG    32'h00000229
`define GTYP_QUAD__CH3_ADAPT_LOP_CFG_SZ 32

`define GTYP_QUAD__CH3_ADAPT_OS_CFG    32'h0000022a
`define GTYP_QUAD__CH3_ADAPT_OS_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_ILO_CFG    32'h0000022b
`define GTYP_QUAD__CH3_CHCLK_ILO_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_MISC_CFG    32'h0000022c
`define GTYP_QUAD__CH3_CHCLK_MISC_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_RSV_CFG    32'h0000022d
`define GTYP_QUAD__CH3_CHCLK_RSV_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG    32'h0000022e
`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG1    32'h0000022f
`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG1_SZ 32

`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG2    32'h00000230
`define GTYP_QUAD__CH3_CHCLK_RXCAL_CFG2_SZ 32

`define GTYP_QUAD__CH3_CHCLK_RXPI_CFG    32'h00000231
`define GTYP_QUAD__CH3_CHCLK_RXPI_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_TXCAL_CFG    32'h00000232
`define GTYP_QUAD__CH3_CHCLK_TXCAL_CFG_SZ 32

`define GTYP_QUAD__CH3_CHCLK_TXPI_CFG0    32'h00000233
`define GTYP_QUAD__CH3_CHCLK_TXPI_CFG0_SZ 32

`define GTYP_QUAD__CH3_CHL_RSV_CFG0    32'h00000234
`define GTYP_QUAD__CH3_CHL_RSV_CFG0_SZ 32

`define GTYP_QUAD__CH3_CHL_RSV_CFG1    32'h00000235
`define GTYP_QUAD__CH3_CHL_RSV_CFG1_SZ 32

`define GTYP_QUAD__CH3_CHL_RSV_CFG2    32'h00000236
`define GTYP_QUAD__CH3_CHL_RSV_CFG2_SZ 32

`define GTYP_QUAD__CH3_CHL_RSV_CFG3    32'h00000237
`define GTYP_QUAD__CH3_CHL_RSV_CFG3_SZ 32

`define GTYP_QUAD__CH3_CHL_RSV_CFG4    32'h00000238
`define GTYP_QUAD__CH3_CHL_RSV_CFG4_SZ 32

`define GTYP_QUAD__CH3_DA_CFG    32'h00000239
`define GTYP_QUAD__CH3_DA_CFG_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG0    32'h0000023a
`define GTYP_QUAD__CH3_EYESCAN_CFG0_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG1    32'h0000023b
`define GTYP_QUAD__CH3_EYESCAN_CFG1_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG10    32'h0000023c
`define GTYP_QUAD__CH3_EYESCAN_CFG10_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG11    32'h0000023d
`define GTYP_QUAD__CH3_EYESCAN_CFG11_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG12    32'h0000023e
`define GTYP_QUAD__CH3_EYESCAN_CFG12_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG13    32'h0000023f
`define GTYP_QUAD__CH3_EYESCAN_CFG13_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG14    32'h00000240
`define GTYP_QUAD__CH3_EYESCAN_CFG14_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG15    32'h00000241
`define GTYP_QUAD__CH3_EYESCAN_CFG15_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG16    32'h00000242
`define GTYP_QUAD__CH3_EYESCAN_CFG16_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG2    32'h00000243
`define GTYP_QUAD__CH3_EYESCAN_CFG2_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG3    32'h00000244
`define GTYP_QUAD__CH3_EYESCAN_CFG3_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG4    32'h00000245
`define GTYP_QUAD__CH3_EYESCAN_CFG4_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG5    32'h00000246
`define GTYP_QUAD__CH3_EYESCAN_CFG5_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG6    32'h00000247
`define GTYP_QUAD__CH3_EYESCAN_CFG6_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG7    32'h00000248
`define GTYP_QUAD__CH3_EYESCAN_CFG7_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG8    32'h00000249
`define GTYP_QUAD__CH3_EYESCAN_CFG8_SZ 32

`define GTYP_QUAD__CH3_EYESCAN_CFG9    32'h0000024a
`define GTYP_QUAD__CH3_EYESCAN_CFG9_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG0    32'h0000024b
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG0_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG1    32'h0000024c
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG1_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG2    32'h0000024d
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG2_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG3    32'h0000024e
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG3_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG4    32'h0000024f
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG4_SZ 32

`define GTYP_QUAD__CH3_FABRIC_INTF_CFG5    32'h00000250
`define GTYP_QUAD__CH3_FABRIC_INTF_CFG5_SZ 32

`define GTYP_QUAD__CH3_INSTANTIATED    32'h00000251
`define GTYP_QUAD__CH3_INSTANTIATED_SZ 1

`define GTYP_QUAD__CH3_MONITOR_CFG    32'h00000252
`define GTYP_QUAD__CH3_MONITOR_CFG_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG0    32'h00000253
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG0_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG1    32'h00000254
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG1_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG10    32'h00000255
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG10_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG2    32'h00000256
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG2_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG3    32'h00000257
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG3_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG4    32'h00000258
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG4_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG5    32'h00000259
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG5_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG6    32'h0000025a
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG6_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG7    32'h0000025b
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG7_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG8    32'h0000025c
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG8_SZ 32

`define GTYP_QUAD__CH3_PIPE_CTRL_CFG9    32'h0000025d
`define GTYP_QUAD__CH3_PIPE_CTRL_CFG9_SZ 32

`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG0    32'h0000025e
`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG0_SZ 32

`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG1    32'h0000025f
`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG1_SZ 32

`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG2    32'h00000260
`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG2_SZ 32

`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG3    32'h00000261
`define GTYP_QUAD__CH3_PIPE_TX_EQ_CFG3_SZ 32

`define GTYP_QUAD__CH3_RESET_BYP_HDSHK_CFG    32'h00000262
`define GTYP_QUAD__CH3_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYP_QUAD__CH3_RESET_CFG    32'h00000263
`define GTYP_QUAD__CH3_RESET_CFG_SZ 32

`define GTYP_QUAD__CH3_RESET_LOOPER_ID_CFG    32'h00000264
`define GTYP_QUAD__CH3_RESET_LOOPER_ID_CFG_SZ 32

`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG0    32'h00000265
`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG0_SZ 32

`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG1    32'h00000266
`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG1_SZ 32

`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG2    32'h00000267
`define GTYP_QUAD__CH3_RESET_LOOP_ID_CFG2_SZ 32

`define GTYP_QUAD__CH3_RESET_TIME_CFG0    32'h00000268
`define GTYP_QUAD__CH3_RESET_TIME_CFG0_SZ 32

`define GTYP_QUAD__CH3_RESET_TIME_CFG1    32'h00000269
`define GTYP_QUAD__CH3_RESET_TIME_CFG1_SZ 32

`define GTYP_QUAD__CH3_RESET_TIME_CFG2    32'h0000026a
`define GTYP_QUAD__CH3_RESET_TIME_CFG2_SZ 32

`define GTYP_QUAD__CH3_RESET_TIME_CFG3    32'h0000026b
`define GTYP_QUAD__CH3_RESET_TIME_CFG3_SZ 32

`define GTYP_QUAD__CH3_RXOUTCLK_FREQ    32'h0000026c
`define GTYP_QUAD__CH3_RXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH3_RXOUTCLK_REF_FREQ    32'h0000026d
`define GTYP_QUAD__CH3_RXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH3_RXOUTCLK_REF_SOURCE    32'h0000026e
`define GTYP_QUAD__CH3_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH3_RX_CDR_CFG0    32'h0000026f
`define GTYP_QUAD__CH3_RX_CDR_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_CDR_CFG1    32'h00000270
`define GTYP_QUAD__CH3_RX_CDR_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_CDR_CFG2    32'h00000271
`define GTYP_QUAD__CH3_RX_CDR_CFG2_SZ 32

`define GTYP_QUAD__CH3_RX_CDR_CFG3    32'h00000272
`define GTYP_QUAD__CH3_RX_CDR_CFG3_SZ 32

`define GTYP_QUAD__CH3_RX_CDR_CFG4    32'h00000273
`define GTYP_QUAD__CH3_RX_CDR_CFG4_SZ 32

`define GTYP_QUAD__CH3_RX_CRC_CFG0    32'h00000274
`define GTYP_QUAD__CH3_RX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_CRC_CFG1    32'h00000275
`define GTYP_QUAD__CH3_RX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_CRC_CFG2    32'h00000276
`define GTYP_QUAD__CH3_RX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH3_RX_CRC_CFG3    32'h00000277
`define GTYP_QUAD__CH3_RX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH3_RX_CTLE_CFG0    32'h00000278
`define GTYP_QUAD__CH3_RX_CTLE_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_CTLE_CFG1    32'h00000279
`define GTYP_QUAD__CH3_RX_CTLE_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_DACI2V_CFG0    32'h0000027a
`define GTYP_QUAD__CH3_RX_DACI2V_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_DATA_RATE    32'h0000027b
`define GTYP_QUAD__CH3_RX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH3_RX_DFE_CFG0    32'h0000027c
`define GTYP_QUAD__CH3_RX_DFE_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG0    32'h0000027d
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG1    32'h0000027e
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG2    32'h0000027f
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG3    32'h00000280
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG4    32'h00000281
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG5    32'h00000282
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG6    32'h00000283
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG7    32'h00000284
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG8    32'h00000285
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG9    32'h00000286
`define GTYP_QUAD__CH3_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYP_QUAD__CH3_RX_MISC_CFG0    32'h00000287
`define GTYP_QUAD__CH3_RX_MISC_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_OOB_CFG0    32'h00000288
`define GTYP_QUAD__CH3_RX_OOB_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_OOB_CFG1    32'h00000289
`define GTYP_QUAD__CH3_RX_OOB_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_PAD_CFG0    32'h0000028a
`define GTYP_QUAD__CH3_RX_PAD_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_PAD_CFG1    32'h0000028b
`define GTYP_QUAD__CH3_RX_PAD_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_PCS_CFG0    32'h0000028c
`define GTYP_QUAD__CH3_RX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_PCS_CFG1    32'h0000028d
`define GTYP_QUAD__CH3_RX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_PCS_CFG2    32'h0000028e
`define GTYP_QUAD__CH3_RX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH3_RX_PCS_CFG3    32'h0000028f
`define GTYP_QUAD__CH3_RX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH3_RX_PCS_CFG4    32'h00000290
`define GTYP_QUAD__CH3_RX_PCS_CFG4_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG0    32'h00000291
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG1    32'h00000292
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG2    32'h00000293
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG3    32'h00000294
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG4    32'h00000295
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH3_RX_PHALIGN_CFG5    32'h00000296
`define GTYP_QUAD__CH3_RX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH3_SIM_MODE    32'h00000297
`define GTYP_QUAD__CH3_SIM_MODE_SZ 48

`define GTYP_QUAD__CH3_SIM_RECEIVER_DETECT_PASS    32'h00000298
`define GTYP_QUAD__CH3_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYP_QUAD__CH3_SIM_RESET_SPEEDUP    32'h00000299
`define GTYP_QUAD__CH3_SIM_RESET_SPEEDUP_SZ 40

`define GTYP_QUAD__CH3_SIM_TX_EIDLE_DRIVE_LEVEL    32'h0000029a
`define GTYP_QUAD__CH3_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYP_QUAD__CH3_TXOUTCLK_FREQ    32'h0000029b
`define GTYP_QUAD__CH3_TXOUTCLK_FREQ_SZ 64

`define GTYP_QUAD__CH3_TXOUTCLK_REF_FREQ    32'h0000029c
`define GTYP_QUAD__CH3_TXOUTCLK_REF_FREQ_SZ 64

`define GTYP_QUAD__CH3_TXOUTCLK_REF_SOURCE    32'h0000029d
`define GTYP_QUAD__CH3_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYP_QUAD__CH3_TX_10G_CFG0    32'h0000029e
`define GTYP_QUAD__CH3_TX_10G_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_10G_CFG1    32'h0000029f
`define GTYP_QUAD__CH3_TX_10G_CFG1_SZ 32

`define GTYP_QUAD__CH3_TX_10G_CFG2    32'h000002a0
`define GTYP_QUAD__CH3_TX_10G_CFG2_SZ 32

`define GTYP_QUAD__CH3_TX_10G_CFG3    32'h000002a1
`define GTYP_QUAD__CH3_TX_10G_CFG3_SZ 32

`define GTYP_QUAD__CH3_TX_ANA_CFG0    32'h000002a2
`define GTYP_QUAD__CH3_TX_ANA_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_CRC_CFG0    32'h000002a3
`define GTYP_QUAD__CH3_TX_CRC_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_CRC_CFG1    32'h000002a4
`define GTYP_QUAD__CH3_TX_CRC_CFG1_SZ 32

`define GTYP_QUAD__CH3_TX_CRC_CFG2    32'h000002a5
`define GTYP_QUAD__CH3_TX_CRC_CFG2_SZ 32

`define GTYP_QUAD__CH3_TX_CRC_CFG3    32'h000002a6
`define GTYP_QUAD__CH3_TX_CRC_CFG3_SZ 32

`define GTYP_QUAD__CH3_TX_DATA_RATE    32'h000002a7
`define GTYP_QUAD__CH3_TX_DATA_RATE_SZ 64

`define GTYP_QUAD__CH3_TX_DRV_CFG0    32'h000002a8
`define GTYP_QUAD__CH3_TX_DRV_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_DRV_CFG1    32'h000002a9
`define GTYP_QUAD__CH3_TX_DRV_CFG1_SZ 32

`define GTYP_QUAD__CH3_TX_PCS_CFG0    32'h000002aa
`define GTYP_QUAD__CH3_TX_PCS_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_PCS_CFG1    32'h000002ab
`define GTYP_QUAD__CH3_TX_PCS_CFG1_SZ 32

`define GTYP_QUAD__CH3_TX_PCS_CFG2    32'h000002ac
`define GTYP_QUAD__CH3_TX_PCS_CFG2_SZ 32

`define GTYP_QUAD__CH3_TX_PCS_CFG3    32'h000002ad
`define GTYP_QUAD__CH3_TX_PCS_CFG3_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG0    32'h000002ae
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG0_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG1    32'h000002af
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG1_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG2    32'h000002b0
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG2_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG3    32'h000002b1
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG3_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG4    32'h000002b2
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG4_SZ 32

`define GTYP_QUAD__CH3_TX_PHALIGN_CFG5    32'h000002b3
`define GTYP_QUAD__CH3_TX_PHALIGN_CFG5_SZ 32

`define GTYP_QUAD__CH3_TX_PIPPM_CFG    32'h000002b4
`define GTYP_QUAD__CH3_TX_PIPPM_CFG_SZ 32

`define GTYP_QUAD__CH3_TX_SER_CFG0    32'h000002b5
`define GTYP_QUAD__CH3_TX_SER_CFG0_SZ 32

`define GTYP_QUAD__CHANNEL_CONNECTIVITY    32'h000002b6
`define GTYP_QUAD__CHANNEL_CONNECTIVITY_SZ 32

`define GTYP_QUAD__CTRL_RSV_CFG0    32'h000002b7
`define GTYP_QUAD__CTRL_RSV_CFG0_SZ 32

`define GTYP_QUAD__CTRL_RSV_CFG1    32'h000002b8
`define GTYP_QUAD__CTRL_RSV_CFG1_SZ 32

`define GTYP_QUAD__HS0_LCPLL_IPS_PIN_EN    32'h000002b9
`define GTYP_QUAD__HS0_LCPLL_IPS_PIN_EN_SZ 1

`define GTYP_QUAD__HS0_LCPLL_IPS_REFCLK_SEL    32'h000002ba
`define GTYP_QUAD__HS0_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP0    32'h000002bb
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP0_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP1    32'h000002bc
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP1_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP2    32'h000002bd
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP2_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP3    32'h000002be
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP3_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP4    32'h000002bf
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP4_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP5    32'h000002c0
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP5_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP6    32'h000002c1
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP6_SZ 3

`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP7    32'h000002c2
`define GTYP_QUAD__HS0_LCPLL_REFCLK_MAP7_SZ 3

`define GTYP_QUAD__HS0_RPLL_IPS_PIN_EN    32'h000002c3
`define GTYP_QUAD__HS0_RPLL_IPS_PIN_EN_SZ 1

`define GTYP_QUAD__HS0_RPLL_IPS_REFCLK_SEL    32'h000002c4
`define GTYP_QUAD__HS0_RPLL_IPS_REFCLK_SEL_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP0    32'h000002c5
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP0_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP1    32'h000002c6
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP1_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP2    32'h000002c7
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP2_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP3    32'h000002c8
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP3_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP4    32'h000002c9
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP4_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP5    32'h000002ca
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP5_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP6    32'h000002cb
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP6_SZ 3

`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP7    32'h000002cc
`define GTYP_QUAD__HS0_RPLL_REFCLK_MAP7_SZ 3

`define GTYP_QUAD__HS1_LCPLL_IPS_PIN_EN    32'h000002cd
`define GTYP_QUAD__HS1_LCPLL_IPS_PIN_EN_SZ 1

`define GTYP_QUAD__HS1_LCPLL_IPS_REFCLK_SEL    32'h000002ce
`define GTYP_QUAD__HS1_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP0    32'h000002cf
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP0_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP1    32'h000002d0
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP1_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP2    32'h000002d1
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP2_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP3    32'h000002d2
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP3_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP4    32'h000002d3
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP4_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP5    32'h000002d4
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP5_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP6    32'h000002d5
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP6_SZ 3

`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP7    32'h000002d6
`define GTYP_QUAD__HS1_LCPLL_REFCLK_MAP7_SZ 3

`define GTYP_QUAD__HS1_RPLL_IPS_PIN_EN    32'h000002d7
`define GTYP_QUAD__HS1_RPLL_IPS_PIN_EN_SZ 1

`define GTYP_QUAD__HS1_RPLL_IPS_REFCLK_SEL    32'h000002d8
`define GTYP_QUAD__HS1_RPLL_IPS_REFCLK_SEL_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP0    32'h000002d9
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP0_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP1    32'h000002da
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP1_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP2    32'h000002db
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP2_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP3    32'h000002dc
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP3_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP4    32'h000002dd
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP4_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP5    32'h000002de
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP5_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP6    32'h000002df
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP6_SZ 3

`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP7    32'h000002e0
`define GTYP_QUAD__HS1_RPLL_REFCLK_MAP7_SZ 3

`define GTYP_QUAD__HSCLK0_HSDIST_CFG    32'h000002e1
`define GTYP_QUAD__HSCLK0_HSDIST_CFG_SZ 32

`define GTYP_QUAD__HSCLK0_INSTANTIATED    32'h000002e2
`define GTYP_QUAD__HSCLK0_INSTANTIATED_SZ 1

`define GTYP_QUAD__HSCLK0_LCPLL_CFG0    32'h000002e3
`define GTYP_QUAD__HSCLK0_LCPLL_CFG0_SZ 32

`define GTYP_QUAD__HSCLK0_LCPLL_CFG1    32'h000002e4
`define GTYP_QUAD__HSCLK0_LCPLL_CFG1_SZ 32

`define GTYP_QUAD__HSCLK0_LCPLL_CFG2    32'h000002e5
`define GTYP_QUAD__HSCLK0_LCPLL_CFG2_SZ 32

`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG0    32'h000002e6
`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG0_SZ 32

`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG1    32'h000002e7
`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG1_SZ 32

`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG2    32'h000002e8
`define GTYP_QUAD__HSCLK0_LCPLL_LGC_CFG2_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_CFG0    32'h000002e9
`define GTYP_QUAD__HSCLK0_RPLL_CFG0_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_CFG1    32'h000002ea
`define GTYP_QUAD__HSCLK0_RPLL_CFG1_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_CFG2    32'h000002eb
`define GTYP_QUAD__HSCLK0_RPLL_CFG2_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG0    32'h000002ec
`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG0_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG1    32'h000002ed
`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG1_SZ 32

`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG2    32'h000002ee
`define GTYP_QUAD__HSCLK0_RPLL_LGC_CFG2_SZ 32

`define GTYP_QUAD__HSCLK0_RXRECCLK_SEL    32'h000002ef
`define GTYP_QUAD__HSCLK0_RXRECCLK_SEL_SZ 2

`define GTYP_QUAD__HSCLK1_HSDIST_CFG    32'h000002f0
`define GTYP_QUAD__HSCLK1_HSDIST_CFG_SZ 32

`define GTYP_QUAD__HSCLK1_INSTANTIATED    32'h000002f1
`define GTYP_QUAD__HSCLK1_INSTANTIATED_SZ 1

`define GTYP_QUAD__HSCLK1_LCPLL_CFG0    32'h000002f2
`define GTYP_QUAD__HSCLK1_LCPLL_CFG0_SZ 32

`define GTYP_QUAD__HSCLK1_LCPLL_CFG1    32'h000002f3
`define GTYP_QUAD__HSCLK1_LCPLL_CFG1_SZ 32

`define GTYP_QUAD__HSCLK1_LCPLL_CFG2    32'h000002f4
`define GTYP_QUAD__HSCLK1_LCPLL_CFG2_SZ 32

`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG0    32'h000002f5
`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG0_SZ 32

`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG1    32'h000002f6
`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG1_SZ 32

`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG2    32'h000002f7
`define GTYP_QUAD__HSCLK1_LCPLL_LGC_CFG2_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_CFG0    32'h000002f8
`define GTYP_QUAD__HSCLK1_RPLL_CFG0_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_CFG1    32'h000002f9
`define GTYP_QUAD__HSCLK1_RPLL_CFG1_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_CFG2    32'h000002fa
`define GTYP_QUAD__HSCLK1_RPLL_CFG2_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG0    32'h000002fb
`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG0_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG1    32'h000002fc
`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG1_SZ 32

`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG2    32'h000002fd
`define GTYP_QUAD__HSCLK1_RPLL_LGC_CFG2_SZ 32

`define GTYP_QUAD__HSCLK1_RXRECCLK_SEL    32'h000002fe
`define GTYP_QUAD__HSCLK1_RXRECCLK_SEL_SZ 2

`define GTYP_QUAD__MEMORY_INIT_FILE    32'h000002ff
`define GTYP_QUAD__MEMORY_INIT_FILE_SZ 32

`define GTYP_QUAD__MST_RESET_CFG    32'h00000300
`define GTYP_QUAD__MST_RESET_CFG_SZ 32

`define GTYP_QUAD__PIN_CFG0    32'h00000301
`define GTYP_QUAD__PIN_CFG0_SZ 32

`define GTYP_QUAD__POR_CFG    32'h00000302
`define GTYP_QUAD__POR_CFG_SZ 32

`define GTYP_QUAD__QUAD_INSTANTIATED    32'h00000303
`define GTYP_QUAD__QUAD_INSTANTIATED_SZ 1

`define GTYP_QUAD__QUAD_SIM_MODE    32'h00000304
`define GTYP_QUAD__QUAD_SIM_MODE_SZ 48

`define GTYP_QUAD__QUAD_SIM_RESET_SPEEDUP    32'h00000305
`define GTYP_QUAD__QUAD_SIM_RESET_SPEEDUP_SZ 40

`define GTYP_QUAD__RCALBG0_CFG0    32'h00000306
`define GTYP_QUAD__RCALBG0_CFG0_SZ 32

`define GTYP_QUAD__RCALBG0_CFG1    32'h00000307
`define GTYP_QUAD__RCALBG0_CFG1_SZ 32

`define GTYP_QUAD__RCALBG0_CFG2    32'h00000308
`define GTYP_QUAD__RCALBG0_CFG2_SZ 32

`define GTYP_QUAD__RCALBG0_CFG3    32'h00000309
`define GTYP_QUAD__RCALBG0_CFG3_SZ 32

`define GTYP_QUAD__RCALBG0_CFG4    32'h0000030a
`define GTYP_QUAD__RCALBG0_CFG4_SZ 32

`define GTYP_QUAD__RCALBG0_CFG5    32'h0000030b
`define GTYP_QUAD__RCALBG0_CFG5_SZ 32

`define GTYP_QUAD__RCALBG1_CFG0    32'h0000030c
`define GTYP_QUAD__RCALBG1_CFG0_SZ 32

`define GTYP_QUAD__RCALBG1_CFG1    32'h0000030d
`define GTYP_QUAD__RCALBG1_CFG1_SZ 32

`define GTYP_QUAD__RCALBG1_CFG2    32'h0000030e
`define GTYP_QUAD__RCALBG1_CFG2_SZ 32

`define GTYP_QUAD__RCALBG1_CFG3    32'h0000030f
`define GTYP_QUAD__RCALBG1_CFG3_SZ 32

`define GTYP_QUAD__RCALBG1_CFG4    32'h00000310
`define GTYP_QUAD__RCALBG1_CFG4_SZ 32

`define GTYP_QUAD__RCALBG1_CFG5    32'h00000311
`define GTYP_QUAD__RCALBG1_CFG5_SZ 32

`define GTYP_QUAD__RXRSTDONE_DIST_SEL    32'h00000312
`define GTYP_QUAD__RXRSTDONE_DIST_SEL_SZ 32

`define GTYP_QUAD__SIM_VERSION    32'h00000313
`define GTYP_QUAD__SIM_VERSION_SZ 2

`define GTYP_QUAD__STAT_NPI_REG_LIST    32'h00000314
`define GTYP_QUAD__STAT_NPI_REG_LIST_SZ 32

`define GTYP_QUAD__TERMPROG_CFG    32'h00000315
`define GTYP_QUAD__TERMPROG_CFG_SZ 32

`define GTYP_QUAD__TXRSTDONE_DIST_SEL    32'h00000316
`define GTYP_QUAD__TXRSTDONE_DIST_SEL_SZ 32

`define GTYP_QUAD__UB_CFG0    32'h00000317
`define GTYP_QUAD__UB_CFG0_SZ 32

`endif  // B_GTYP_QUAD_DEFINES_VH