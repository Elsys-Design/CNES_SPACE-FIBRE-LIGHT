// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     blh_composer 3.0001
//    Built On:     Tue Aug 30 09:51:45 2016
//    Bundle:       PCIE40E4
//    Architecture: diablo
//    Snapshot Dir: /tmp/mu8kpKnzTO
// Environment Variables:
//    XILENV=""
//    MYXILENV=""
//

`ifdef B_PCIE40E4_DEFINES_VH
`else
`define B_PCIE40E4_DEFINES_VH

// Look-up table parameters
//

`define PCIE40E4_ADDR_N  520
`define PCIE40E4_ADDR_SZ 32
`define PCIE40E4_DATA_SZ 152

// Attribute addresses
//

`define PCIE40E4__ARI_CAP_ENABLE   	32'h0000	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__ARI_CAP_ENABLE_SZ	40

`define PCIE40E4__AUTO_FLR_RESPONSE   	32'h0001	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AUTO_FLR_RESPONSE_SZ	40

`define PCIE40E4__AXISTEN_IF_CC_ALIGNMENT_MODE   	32'h0002	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__AXISTEN_IF_CC_ALIGNMENT_MODE_SZ	2

`define PCIE40E4__AXISTEN_IF_COMPL_TIMEOUT_REG0   	32'h0003	// Type=HEX; Min=24'h000000, Max=24'hffffff
`define PCIE40E4__AXISTEN_IF_COMPL_TIMEOUT_REG0_SZ	24

`define PCIE40E4__AXISTEN_IF_COMPL_TIMEOUT_REG1   	32'h0004	// Type=HEX; Min=28'h0000000, Max=28'hfffffff
`define PCIE40E4__AXISTEN_IF_COMPL_TIMEOUT_REG1_SZ	28

`define PCIE40E4__AXISTEN_IF_CQ_ALIGNMENT_MODE   	32'h0005	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__AXISTEN_IF_CQ_ALIGNMENT_MODE_SZ	2

`define PCIE40E4__AXISTEN_IF_CQ_EN_POISONED_MEM_WR   	32'h0006	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_CQ_EN_POISONED_MEM_WR_SZ	40

`define PCIE40E4__AXISTEN_IF_ENABLE_256_TAGS   	32'h0007	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_ENABLE_256_TAGS_SZ	40

`define PCIE40E4__AXISTEN_IF_ENABLE_CLIENT_TAG   	32'h0008	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_ENABLE_CLIENT_TAG_SZ	40

`define PCIE40E4__AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE   	32'h0009	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE_SZ	40

`define PCIE40E4__AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK   	32'h000a	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK_SZ	40

`define PCIE40E4__AXISTEN_IF_ENABLE_MSG_ROUTE   	32'h000b	// Type=HEX; Min=18'h00000, Max=18'h3ffff
`define PCIE40E4__AXISTEN_IF_ENABLE_MSG_ROUTE_SZ	18

`define PCIE40E4__AXISTEN_IF_ENABLE_RX_MSG_INTFC   	32'h000c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_ENABLE_RX_MSG_INTFC_SZ	40

`define PCIE40E4__AXISTEN_IF_EXT_512   	32'h000d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_EXT_512_SZ	40

`define PCIE40E4__AXISTEN_IF_EXT_512_CC_STRADDLE   	32'h000e	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_EXT_512_CC_STRADDLE_SZ	40

`define PCIE40E4__AXISTEN_IF_EXT_512_CQ_STRADDLE   	32'h000f	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_EXT_512_CQ_STRADDLE_SZ	40

`define PCIE40E4__AXISTEN_IF_EXT_512_RC_STRADDLE   	32'h0010	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_EXT_512_RC_STRADDLE_SZ	40

`define PCIE40E4__AXISTEN_IF_EXT_512_RQ_STRADDLE   	32'h0011	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_EXT_512_RQ_STRADDLE_SZ	40

`define PCIE40E4__AXISTEN_IF_LEGACY_MODE_ENABLE   	32'h0012	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_LEGACY_MODE_ENABLE_SZ	40

`define PCIE40E4__AXISTEN_IF_MSIX_FROM_RAM_PIPELINE   	32'h0013	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_MSIX_FROM_RAM_PIPELINE_SZ	40

`define PCIE40E4__AXISTEN_IF_MSIX_RX_PARITY_EN   	32'h0014	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__AXISTEN_IF_MSIX_RX_PARITY_EN_SZ	40

`define PCIE40E4__AXISTEN_IF_MSIX_TO_RAM_PIPELINE   	32'h0015	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_MSIX_TO_RAM_PIPELINE_SZ	40

`define PCIE40E4__AXISTEN_IF_RC_ALIGNMENT_MODE   	32'h0016	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__AXISTEN_IF_RC_ALIGNMENT_MODE_SZ	2

`define PCIE40E4__AXISTEN_IF_RC_STRADDLE   	32'h0017	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_RC_STRADDLE_SZ	40

`define PCIE40E4__AXISTEN_IF_RQ_ALIGNMENT_MODE   	32'h0018	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__AXISTEN_IF_RQ_ALIGNMENT_MODE_SZ	2

`define PCIE40E4__AXISTEN_IF_RX_PARITY_EN   	32'h0019	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__AXISTEN_IF_RX_PARITY_EN_SZ	40

`define PCIE40E4__AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT   	32'h001a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT_SZ	40

`define PCIE40E4__AXISTEN_IF_TX_PARITY_EN   	32'h001b	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__AXISTEN_IF_TX_PARITY_EN_SZ	40

`define PCIE40E4__AXISTEN_IF_WIDTH   	32'h001c	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__AXISTEN_IF_WIDTH_SZ	2

`define PCIE40E4__CFG_BYPASS_MODE_ENABLE   	32'h001d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__CFG_BYPASS_MODE_ENABLE_SZ	40

`define PCIE40E4__CRM_CORE_CLK_FREQ_500   	32'h001e	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__CRM_CORE_CLK_FREQ_500_SZ	40

`define PCIE40E4__CRM_USER_CLK_FREQ   	32'h001f	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__CRM_USER_CLK_FREQ_SZ	2

`define PCIE40E4__DEBUG_AXI4ST_SPARE   	32'h0020	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__DEBUG_AXI4ST_SPARE_SZ	16

`define PCIE40E4__DEBUG_AXIST_DISABLE_FEATURE_BIT   	32'h0021	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__DEBUG_AXIST_DISABLE_FEATURE_BIT_SZ	8

`define PCIE40E4__DEBUG_CAR_SPARE   	32'h0022	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__DEBUG_CAR_SPARE_SZ	4

`define PCIE40E4__DEBUG_CFG_SPARE   	32'h0023	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__DEBUG_CFG_SPARE_SZ	16

`define PCIE40E4__DEBUG_LL_SPARE   	32'h0024	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__DEBUG_LL_SPARE_SZ	16

`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR   	32'h0025	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR_SZ	40

`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR   	32'h0026	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR_SZ	40

`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR   	32'h0027	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR_SZ	40

`define PCIE40E4__DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL   	32'h0028	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL_SZ	40

`define PCIE40E4__DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW   	32'h0029	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW_SZ	40

`define PCIE40E4__DEBUG_PL_DISABLE_SCRAMBLING   	32'h002a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_DISABLE_SCRAMBLING_SZ	40

`define PCIE40E4__DEBUG_PL_SIM_RESET_LFSR   	32'h002b	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_PL_SIM_RESET_LFSR_SZ	40

`define PCIE40E4__DEBUG_PL_SPARE   	32'h002c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__DEBUG_PL_SPARE_SZ	16

`define PCIE40E4__DEBUG_TL_DISABLE_FC_TIMEOUT   	32'h002d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_TL_DISABLE_FC_TIMEOUT_SZ	40

`define PCIE40E4__DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS   	32'h002e	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_SZ	40

`define PCIE40E4__DEBUG_TL_SPARE   	32'h002f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__DEBUG_TL_SPARE_SZ	16

`define PCIE40E4__DNSTREAM_LINK_NUM   	32'h0030	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__DNSTREAM_LINK_NUM_SZ	8

`define PCIE40E4__DSN_CAP_ENABLE   	32'h0031	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__DSN_CAP_ENABLE_SZ	40

`define PCIE40E4__EXTENDED_CFG_EXTEND_INTERFACE_ENABLE   	32'h0032	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_SZ	40

`define PCIE40E4__HEADER_TYPE_OVERRIDE   	32'h0033	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__HEADER_TYPE_OVERRIDE_SZ	40

`define PCIE40E4__IS_SWITCH_PORT   	32'h0034	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__IS_SWITCH_PORT_SZ	40

`define PCIE40E4__LEGACY_CFG_EXTEND_INTERFACE_ENABLE   	32'h0035	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LEGACY_CFG_EXTEND_INTERFACE_ENABLE_SZ	40

`define PCIE40E4__LL_ACK_TIMEOUT   	32'h0036	// Type=HEX; Min=9'h000, Max=9'h1ff
`define PCIE40E4__LL_ACK_TIMEOUT_SZ	9

`define PCIE40E4__LL_ACK_TIMEOUT_EN   	32'h0037	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LL_ACK_TIMEOUT_EN_SZ	40

`define PCIE40E4__LL_ACK_TIMEOUT_FUNC   	32'h0038	// Type=DECIMAL; Values=0,1,2,3
`define PCIE40E4__LL_ACK_TIMEOUT_FUNC_SZ	32

`define PCIE40E4__LL_DISABLE_SCHED_TX_NAK   	32'h0039	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LL_DISABLE_SCHED_TX_NAK_SZ	40

`define PCIE40E4__LL_REPLAY_FROM_RAM_PIPELINE   	32'h003a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LL_REPLAY_FROM_RAM_PIPELINE_SZ	40

`define PCIE40E4__LL_REPLAY_TIMEOUT   	32'h003b	// Type=HEX; Min=9'h000, Max=9'h1ff
`define PCIE40E4__LL_REPLAY_TIMEOUT_SZ	9

`define PCIE40E4__LL_REPLAY_TIMEOUT_EN   	32'h003c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LL_REPLAY_TIMEOUT_EN_SZ	40

`define PCIE40E4__LL_REPLAY_TIMEOUT_FUNC   	32'h003d	// Type=DECIMAL; Values=0,1,2,3
`define PCIE40E4__LL_REPLAY_TIMEOUT_FUNC_SZ	32

`define PCIE40E4__LL_REPLAY_TO_RAM_PIPELINE   	32'h003e	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LL_REPLAY_TO_RAM_PIPELINE_SZ	40

`define PCIE40E4__LL_RX_TLP_PARITY_GEN   	32'h003f	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__LL_RX_TLP_PARITY_GEN_SZ	40

`define PCIE40E4__LL_TX_TLP_PARITY_CHK   	32'h0040	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__LL_TX_TLP_PARITY_CHK_SZ	40

`define PCIE40E4__LL_USER_SPARE   	32'h0041	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__LL_USER_SPARE_SZ	16

`define PCIE40E4__LTR_TX_MESSAGE_MINIMUM_INTERVAL   	32'h0042	// Type=HEX; Min=10'h000, Max=10'h3ff
`define PCIE40E4__LTR_TX_MESSAGE_MINIMUM_INTERVAL_SZ	10

`define PCIE40E4__LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE   	32'h0043	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_SZ	40

`define PCIE40E4__LTR_TX_MESSAGE_ON_LTR_ENABLE   	32'h0044	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__LTR_TX_MESSAGE_ON_LTR_ENABLE_SZ	40

`define PCIE40E4__MCAP_CAP_NEXTPTR   	32'h0045	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__MCAP_CAP_NEXTPTR_SZ	12

`define PCIE40E4__MCAP_CONFIGURE_OVERRIDE   	32'h0046	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_CONFIGURE_OVERRIDE_SZ	40

`define PCIE40E4__MCAP_ENABLE   	32'h0047	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_ENABLE_SZ	40

`define PCIE40E4__MCAP_EOS_DESIGN_SWITCH   	32'h0048	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_EOS_DESIGN_SWITCH_SZ	40

`define PCIE40E4__MCAP_FPGA_BITSTREAM_VERSION   	32'h0049	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__MCAP_FPGA_BITSTREAM_VERSION_SZ	32

`define PCIE40E4__MCAP_GATE_IO_ENABLE_DESIGN_SWITCH   	32'h004a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_SZ	40

`define PCIE40E4__MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH   	32'h004b	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_SZ	40

`define PCIE40E4__MCAP_INPUT_GATE_DESIGN_SWITCH   	32'h004c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_INPUT_GATE_DESIGN_SWITCH_SZ	40

`define PCIE40E4__MCAP_INTERRUPT_ON_MCAP_EOS   	32'h004d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_INTERRUPT_ON_MCAP_EOS_SZ	40

`define PCIE40E4__MCAP_INTERRUPT_ON_MCAP_ERROR   	32'h004e	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__MCAP_INTERRUPT_ON_MCAP_ERROR_SZ	40

`define PCIE40E4__MCAP_VSEC_ID   	32'h004f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__MCAP_VSEC_ID_SZ	16

`define PCIE40E4__MCAP_VSEC_LEN   	32'h0050	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__MCAP_VSEC_LEN_SZ	12

`define PCIE40E4__MCAP_VSEC_REV   	32'h0051	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__MCAP_VSEC_REV_SZ	4

`define PCIE40E4__PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE   	32'h0052	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE_SZ	40

`define PCIE40E4__PF0_AER_CAP_NEXTPTR   	32'h0053	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_AER_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_ARI_CAP_NEXTPTR   	32'h0054	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_ARI_CAP_NEXT_FUNC   	32'h0055	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_ARI_CAP_NEXT_FUNC_SZ	8

`define PCIE40E4__PF0_ARI_CAP_VER   	32'h0056	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF0_ARI_CAP_VER_SZ	4

`define PCIE40E4__PF0_BAR0_APERTURE_SIZE   	32'h0057	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_BAR0_CONTROL   	32'h0058	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF0_BAR1_APERTURE_SIZE   	32'h0059	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_BAR1_CONTROL   	32'h005a	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF0_BAR2_APERTURE_SIZE   	32'h005b	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_BAR2_CONTROL   	32'h005c	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF0_BAR3_APERTURE_SIZE   	32'h005d	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_BAR3_CONTROL   	32'h005e	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF0_BAR4_APERTURE_SIZE   	32'h005f	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_BAR4_CONTROL   	32'h0060	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF0_BAR5_APERTURE_SIZE   	32'h0061	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_BAR5_CONTROL   	32'h0062	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF0_CAPABILITY_POINTER   	32'h0063	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_CAPABILITY_POINTER_SZ	8

`define PCIE40E4__PF0_CLASS_CODE   	32'h0064	// Type=HEX; Min=24'h000000, Max=24'hffffff
`define PCIE40E4__PF0_CLASS_CODE_SZ	24

`define PCIE40E4__PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT   	32'h0065	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT   	32'h0066	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT   	32'h0067	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_ARI_FORWARD_ENABLE   	32'h0068	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_DEV_CAP2_ARI_FORWARD_ENABLE_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE   	32'h0069	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_LTR_SUPPORT   	32'h006a	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP2_LTR_SUPPORT_SZ	40

`define PCIE40E4__PF0_DEV_CAP2_OBFF_SUPPORT   	32'h006b	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PF0_DEV_CAP2_OBFF_SUPPORT_SZ	2

`define PCIE40E4__PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT   	32'h006c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_SZ	40

`define PCIE40E4__PF0_DEV_CAP_ENDPOINT_L0S_LATENCY   	32'h006d	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_SZ	32

`define PCIE40E4__PF0_DEV_CAP_ENDPOINT_L1_LATENCY   	32'h006e	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF0_DEV_CAP_ENDPOINT_L1_LATENCY_SZ	32

`define PCIE40E4__PF0_DEV_CAP_EXT_TAG_SUPPORTED   	32'h006f	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP_EXT_TAG_SUPPORTED_SZ	40

`define PCIE40E4__PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE   	32'h0070	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_SZ	40

`define PCIE40E4__PF0_DEV_CAP_MAX_PAYLOAD_SIZE   	32'h0071	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_DEV_CAP_MAX_PAYLOAD_SIZE_SZ	3

`define PCIE40E4__PF0_DSN_CAP_NEXTPTR   	32'h0072	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_DSN_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_EXPANSION_ROM_APERTURE_SIZE   	32'h0073	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_EXPANSION_ROM_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_EXPANSION_ROM_ENABLE   	32'h0074	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_EXPANSION_ROM_ENABLE_SZ	40

`define PCIE40E4__PF0_INTERRUPT_PIN   	32'h0075	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_INTERRUPT_PIN_SZ	3

`define PCIE40E4__PF0_LINK_CAP_ASPM_SUPPORT   	32'h0076	// Type=DECIMAL; Values=0,1,2,3
`define PCIE40E4__PF0_LINK_CAP_ASPM_SUPPORT_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1   	32'h0077	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2   	32'h0078	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3   	32'h0079	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4   	32'h007a	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1   	32'h007b	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2   	32'h007c	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3   	32'h007d	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4   	32'h007e	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1   	32'h007f	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2   	32'h0080	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3   	32'h0081	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4   	32'h0082	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1   	32'h0083	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2   	32'h0084	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3   	32'h0085	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_SZ	32

`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4   	32'h0086	// Type=DECIMAL; Values=7,0,1,2,3,4,5,6
`define PCIE40E4__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4_SZ	32

`define PCIE40E4__PF0_LINK_CONTROL_RCB   	32'h0087	// Type=HEX; Min=1'h0, Max=1'h1
`define PCIE40E4__PF0_LINK_CONTROL_RCB_SZ	1

`define PCIE40E4__PF0_LINK_STATUS_SLOT_CLOCK_CONFIG   	32'h0088	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_SZ	40

`define PCIE40E4__PF0_LTR_CAP_MAX_NOSNOOP_LAT   	32'h0089	// Type=HEX; Min=10'h000, Max=10'h3ff
`define PCIE40E4__PF0_LTR_CAP_MAX_NOSNOOP_LAT_SZ	10

`define PCIE40E4__PF0_LTR_CAP_MAX_SNOOP_LAT   	32'h008a	// Type=HEX; Min=10'h000, Max=10'h3ff
`define PCIE40E4__PF0_LTR_CAP_MAX_SNOOP_LAT_SZ	10

`define PCIE40E4__PF0_LTR_CAP_NEXTPTR   	32'h008b	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_LTR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_LTR_CAP_VER   	32'h008c	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF0_LTR_CAP_VER_SZ	4

`define PCIE40E4__PF0_MSIX_CAP_NEXTPTR   	32'h008d	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF0_MSIX_CAP_PBA_BIR   	32'h008e	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF0_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__PF0_MSIX_CAP_PBA_OFFSET   	32'h008f	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF0_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__PF0_MSIX_CAP_TABLE_BIR   	32'h0090	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF0_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__PF0_MSIX_CAP_TABLE_OFFSET   	32'h0091	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF0_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__PF0_MSIX_CAP_TABLE_SIZE   	32'h0092	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__PF0_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__PF0_MSIX_VECTOR_COUNT   	32'h0093	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_MSIX_VECTOR_COUNT_SZ	6

`define PCIE40E4__PF0_MSI_CAP_MULTIMSGCAP   	32'h0094	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF0_MSI_CAP_MULTIMSGCAP_SZ	32

`define PCIE40E4__PF0_MSI_CAP_NEXTPTR   	32'h0095	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_MSI_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF0_MSI_CAP_PERVECMASKCAP   	32'h0096	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_MSI_CAP_PERVECMASKCAP_SZ	40

`define PCIE40E4__PF0_PCIE_CAP_NEXTPTR   	32'h0097	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF0_PM_CAP_ID   	32'h0098	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_PM_CAP_ID_SZ	8

`define PCIE40E4__PF0_PM_CAP_NEXTPTR   	32'h0099	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF0_PM_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D0   	32'h009a	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D0_SZ	40

`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D1   	32'h009b	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D1_SZ	40

`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D3HOT   	32'h009c	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_PM_CAP_PMESUPPORT_D3HOT_SZ	40

`define PCIE40E4__PF0_PM_CAP_SUPP_D1_STATE   	32'h009d	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_PM_CAP_SUPP_D1_STATE_SZ	40

`define PCIE40E4__PF0_PM_CAP_VER_ID   	32'h009e	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_PM_CAP_VER_ID_SZ	3

`define PCIE40E4__PF0_PM_CSR_NOSOFTRESET   	32'h009f	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_PM_CSR_NOSOFTRESET_SZ	40

`define PCIE40E4__PF0_SECONDARY_PCIE_CAP_NEXTPTR   	32'h00a0	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_SECONDARY_PCIE_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED   	32'h00a1	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ	40

`define PCIE40E4__PF0_SRIOV_BAR0_APERTURE_SIZE   	32'h00a2	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_SRIOV_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_SRIOV_BAR0_CONTROL   	32'h00a3	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_BAR1_APERTURE_SIZE   	32'h00a4	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_SRIOV_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_SRIOV_BAR1_CONTROL   	32'h00a5	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_BAR2_APERTURE_SIZE   	32'h00a6	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_SRIOV_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_SRIOV_BAR2_CONTROL   	32'h00a7	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_BAR3_APERTURE_SIZE   	32'h00a8	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_SRIOV_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_SRIOV_BAR3_CONTROL   	32'h00a9	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_BAR4_APERTURE_SIZE   	32'h00aa	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF0_SRIOV_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF0_SRIOV_BAR4_CONTROL   	32'h00ab	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_BAR5_APERTURE_SIZE   	32'h00ac	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF0_SRIOV_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF0_SRIOV_BAR5_CONTROL   	32'h00ad	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_SRIOV_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF0_SRIOV_CAP_INITIAL_VF   	32'h00ae	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF0_SRIOV_CAP_INITIAL_VF_SZ	16

`define PCIE40E4__PF0_SRIOV_CAP_NEXTPTR   	32'h00af	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_SRIOV_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_SRIOV_CAP_TOTAL_VF   	32'h00b0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF0_SRIOV_CAP_TOTAL_VF_SZ	16

`define PCIE40E4__PF0_SRIOV_CAP_VER   	32'h00b1	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF0_SRIOV_CAP_VER_SZ	4

`define PCIE40E4__PF0_SRIOV_FIRST_VF_OFFSET   	32'h00b2	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF0_SRIOV_FIRST_VF_OFFSET_SZ	16

`define PCIE40E4__PF0_SRIOV_FUNC_DEP_LINK   	32'h00b3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF0_SRIOV_FUNC_DEP_LINK_SZ	16

`define PCIE40E4__PF0_SRIOV_SUPPORTED_PAGE_SIZE   	32'h00b4	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PF0_SRIOV_SUPPORTED_PAGE_SIZE_SZ	32

`define PCIE40E4__PF0_SRIOV_VF_DEVICE_ID   	32'h00b5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF0_SRIOV_VF_DEVICE_ID_SZ	16

`define PCIE40E4__PF0_TPHR_CAP_DEV_SPECIFIC_MODE   	32'h00b6	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_TPHR_CAP_DEV_SPECIFIC_MODE_SZ	40

`define PCIE40E4__PF0_TPHR_CAP_ENABLE   	32'h00b7	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_TPHR_CAP_ENABLE_SZ	40

`define PCIE40E4__PF0_TPHR_CAP_INT_VEC_MODE   	32'h00b8	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PF0_TPHR_CAP_INT_VEC_MODE_SZ	40

`define PCIE40E4__PF0_TPHR_CAP_NEXTPTR   	32'h00b9	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_TPHR_CAP_ST_MODE_SEL   	32'h00ba	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF0_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__PF0_TPHR_CAP_ST_TABLE_LOC   	32'h00bb	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PF0_TPHR_CAP_ST_TABLE_LOC_SZ	2

`define PCIE40E4__PF0_TPHR_CAP_ST_TABLE_SIZE   	32'h00bc	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__PF0_TPHR_CAP_ST_TABLE_SIZE_SZ	11

`define PCIE40E4__PF0_TPHR_CAP_VER   	32'h00bd	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF0_TPHR_CAP_VER_SZ	4

`define PCIE40E4__PF0_VC_CAP_ENABLE   	32'h00be	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF0_VC_CAP_ENABLE_SZ	40

`define PCIE40E4__PF0_VC_CAP_NEXTPTR   	32'h00bf	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF0_VC_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF0_VC_CAP_VER   	32'h00c0	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF0_VC_CAP_VER_SZ	4

`define PCIE40E4__PF1_AER_CAP_NEXTPTR   	32'h00c1	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF1_AER_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF1_ARI_CAP_NEXTPTR   	32'h00c2	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF1_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF1_ARI_CAP_NEXT_FUNC   	32'h00c3	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_ARI_CAP_NEXT_FUNC_SZ	8

`define PCIE40E4__PF1_BAR0_APERTURE_SIZE   	32'h00c4	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_BAR0_CONTROL   	32'h00c5	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF1_BAR1_APERTURE_SIZE   	32'h00c6	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_BAR1_CONTROL   	32'h00c7	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF1_BAR2_APERTURE_SIZE   	32'h00c8	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_BAR2_CONTROL   	32'h00c9	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF1_BAR3_APERTURE_SIZE   	32'h00ca	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_BAR3_CONTROL   	32'h00cb	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF1_BAR4_APERTURE_SIZE   	32'h00cc	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_BAR4_CONTROL   	32'h00cd	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF1_BAR5_APERTURE_SIZE   	32'h00ce	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_BAR5_CONTROL   	32'h00cf	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF1_CAPABILITY_POINTER   	32'h00d0	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_CAPABILITY_POINTER_SZ	8

`define PCIE40E4__PF1_CLASS_CODE   	32'h00d1	// Type=HEX; Min=24'h000000, Max=24'hffffff
`define PCIE40E4__PF1_CLASS_CODE_SZ	24

`define PCIE40E4__PF1_DEV_CAP_MAX_PAYLOAD_SIZE   	32'h00d2	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_DEV_CAP_MAX_PAYLOAD_SIZE_SZ	3

`define PCIE40E4__PF1_DSN_CAP_NEXTPTR   	32'h00d3	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF1_DSN_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF1_EXPANSION_ROM_APERTURE_SIZE   	32'h00d4	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_EXPANSION_ROM_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_EXPANSION_ROM_ENABLE   	32'h00d5	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF1_EXPANSION_ROM_ENABLE_SZ	40

`define PCIE40E4__PF1_INTERRUPT_PIN   	32'h00d6	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_INTERRUPT_PIN_SZ	3

`define PCIE40E4__PF1_MSIX_CAP_NEXTPTR   	32'h00d7	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF1_MSIX_CAP_PBA_BIR   	32'h00d8	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF1_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__PF1_MSIX_CAP_PBA_OFFSET   	32'h00d9	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF1_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__PF1_MSIX_CAP_TABLE_BIR   	32'h00da	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF1_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__PF1_MSIX_CAP_TABLE_OFFSET   	32'h00db	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF1_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__PF1_MSIX_CAP_TABLE_SIZE   	32'h00dc	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__PF1_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__PF1_MSI_CAP_MULTIMSGCAP   	32'h00dd	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF1_MSI_CAP_MULTIMSGCAP_SZ	32

`define PCIE40E4__PF1_MSI_CAP_NEXTPTR   	32'h00de	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_MSI_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF1_MSI_CAP_PERVECMASKCAP   	32'h00df	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF1_MSI_CAP_PERVECMASKCAP_SZ	40

`define PCIE40E4__PF1_PCIE_CAP_NEXTPTR   	32'h00e0	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF1_PM_CAP_NEXTPTR   	32'h00e1	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF1_PM_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED   	32'h00e2	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ	40

`define PCIE40E4__PF1_SRIOV_BAR0_APERTURE_SIZE   	32'h00e3	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_SRIOV_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_SRIOV_BAR0_CONTROL   	32'h00e4	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_BAR1_APERTURE_SIZE   	32'h00e5	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_SRIOV_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_SRIOV_BAR1_CONTROL   	32'h00e6	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_BAR2_APERTURE_SIZE   	32'h00e7	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_SRIOV_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_SRIOV_BAR2_CONTROL   	32'h00e8	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_BAR3_APERTURE_SIZE   	32'h00e9	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_SRIOV_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_SRIOV_BAR3_CONTROL   	32'h00ea	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_BAR4_APERTURE_SIZE   	32'h00eb	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF1_SRIOV_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF1_SRIOV_BAR4_CONTROL   	32'h00ec	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_BAR5_APERTURE_SIZE   	32'h00ed	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF1_SRIOV_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF1_SRIOV_BAR5_CONTROL   	32'h00ee	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_SRIOV_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF1_SRIOV_CAP_INITIAL_VF   	32'h00ef	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF1_SRIOV_CAP_INITIAL_VF_SZ	16

`define PCIE40E4__PF1_SRIOV_CAP_NEXTPTR   	32'h00f0	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF1_SRIOV_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF1_SRIOV_CAP_TOTAL_VF   	32'h00f1	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF1_SRIOV_CAP_TOTAL_VF_SZ	16

`define PCIE40E4__PF1_SRIOV_CAP_VER   	32'h00f2	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF1_SRIOV_CAP_VER_SZ	4

`define PCIE40E4__PF1_SRIOV_FIRST_VF_OFFSET   	32'h00f3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF1_SRIOV_FIRST_VF_OFFSET_SZ	16

`define PCIE40E4__PF1_SRIOV_FUNC_DEP_LINK   	32'h00f4	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF1_SRIOV_FUNC_DEP_LINK_SZ	16

`define PCIE40E4__PF1_SRIOV_SUPPORTED_PAGE_SIZE   	32'h00f5	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PF1_SRIOV_SUPPORTED_PAGE_SIZE_SZ	32

`define PCIE40E4__PF1_SRIOV_VF_DEVICE_ID   	32'h00f6	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF1_SRIOV_VF_DEVICE_ID_SZ	16

`define PCIE40E4__PF1_TPHR_CAP_NEXTPTR   	32'h00f7	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF1_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF1_TPHR_CAP_ST_MODE_SEL   	32'h00f8	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF1_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__PF2_AER_CAP_NEXTPTR   	32'h00f9	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF2_AER_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF2_ARI_CAP_NEXTPTR   	32'h00fa	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF2_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF2_ARI_CAP_NEXT_FUNC   	32'h00fb	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_ARI_CAP_NEXT_FUNC_SZ	8

`define PCIE40E4__PF2_BAR0_APERTURE_SIZE   	32'h00fc	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_BAR0_CONTROL   	32'h00fd	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF2_BAR1_APERTURE_SIZE   	32'h00fe	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_BAR1_CONTROL   	32'h00ff	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF2_BAR2_APERTURE_SIZE   	32'h0100	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_BAR2_CONTROL   	32'h0101	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF2_BAR3_APERTURE_SIZE   	32'h0102	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_BAR3_CONTROL   	32'h0103	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF2_BAR4_APERTURE_SIZE   	32'h0104	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_BAR4_CONTROL   	32'h0105	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF2_BAR5_APERTURE_SIZE   	32'h0106	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_BAR5_CONTROL   	32'h0107	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF2_CAPABILITY_POINTER   	32'h0108	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_CAPABILITY_POINTER_SZ	8

`define PCIE40E4__PF2_CLASS_CODE   	32'h0109	// Type=HEX; Min=24'h000000, Max=24'hffffff
`define PCIE40E4__PF2_CLASS_CODE_SZ	24

`define PCIE40E4__PF2_DEV_CAP_MAX_PAYLOAD_SIZE   	32'h010a	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_DEV_CAP_MAX_PAYLOAD_SIZE_SZ	3

`define PCIE40E4__PF2_DSN_CAP_NEXTPTR   	32'h010b	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF2_DSN_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF2_EXPANSION_ROM_APERTURE_SIZE   	32'h010c	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_EXPANSION_ROM_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_EXPANSION_ROM_ENABLE   	32'h010d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF2_EXPANSION_ROM_ENABLE_SZ	40

`define PCIE40E4__PF2_INTERRUPT_PIN   	32'h010e	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_INTERRUPT_PIN_SZ	3

`define PCIE40E4__PF2_MSIX_CAP_NEXTPTR   	32'h010f	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF2_MSIX_CAP_PBA_BIR   	32'h0110	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF2_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__PF2_MSIX_CAP_PBA_OFFSET   	32'h0111	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF2_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__PF2_MSIX_CAP_TABLE_BIR   	32'h0112	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF2_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__PF2_MSIX_CAP_TABLE_OFFSET   	32'h0113	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF2_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__PF2_MSIX_CAP_TABLE_SIZE   	32'h0114	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__PF2_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__PF2_MSI_CAP_MULTIMSGCAP   	32'h0115	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF2_MSI_CAP_MULTIMSGCAP_SZ	32

`define PCIE40E4__PF2_MSI_CAP_NEXTPTR   	32'h0116	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_MSI_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF2_MSI_CAP_PERVECMASKCAP   	32'h0117	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF2_MSI_CAP_PERVECMASKCAP_SZ	40

`define PCIE40E4__PF2_PCIE_CAP_NEXTPTR   	32'h0118	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF2_PM_CAP_NEXTPTR   	32'h0119	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF2_PM_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED   	32'h011a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ	40

`define PCIE40E4__PF2_SRIOV_BAR0_APERTURE_SIZE   	32'h011b	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_SRIOV_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_SRIOV_BAR0_CONTROL   	32'h011c	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_BAR1_APERTURE_SIZE   	32'h011d	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_SRIOV_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_SRIOV_BAR1_CONTROL   	32'h011e	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_BAR2_APERTURE_SIZE   	32'h011f	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_SRIOV_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_SRIOV_BAR2_CONTROL   	32'h0120	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_BAR3_APERTURE_SIZE   	32'h0121	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_SRIOV_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_SRIOV_BAR3_CONTROL   	32'h0122	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_BAR4_APERTURE_SIZE   	32'h0123	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF2_SRIOV_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF2_SRIOV_BAR4_CONTROL   	32'h0124	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_BAR5_APERTURE_SIZE   	32'h0125	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF2_SRIOV_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF2_SRIOV_BAR5_CONTROL   	32'h0126	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_SRIOV_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF2_SRIOV_CAP_INITIAL_VF   	32'h0127	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF2_SRIOV_CAP_INITIAL_VF_SZ	16

`define PCIE40E4__PF2_SRIOV_CAP_NEXTPTR   	32'h0128	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF2_SRIOV_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF2_SRIOV_CAP_TOTAL_VF   	32'h0129	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF2_SRIOV_CAP_TOTAL_VF_SZ	16

`define PCIE40E4__PF2_SRIOV_CAP_VER   	32'h012a	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF2_SRIOV_CAP_VER_SZ	4

`define PCIE40E4__PF2_SRIOV_FIRST_VF_OFFSET   	32'h012b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF2_SRIOV_FIRST_VF_OFFSET_SZ	16

`define PCIE40E4__PF2_SRIOV_FUNC_DEP_LINK   	32'h012c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF2_SRIOV_FUNC_DEP_LINK_SZ	16

`define PCIE40E4__PF2_SRIOV_SUPPORTED_PAGE_SIZE   	32'h012d	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PF2_SRIOV_SUPPORTED_PAGE_SIZE_SZ	32

`define PCIE40E4__PF2_SRIOV_VF_DEVICE_ID   	32'h012e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF2_SRIOV_VF_DEVICE_ID_SZ	16

`define PCIE40E4__PF2_TPHR_CAP_NEXTPTR   	32'h012f	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF2_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF2_TPHR_CAP_ST_MODE_SEL   	32'h0130	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF2_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__PF3_AER_CAP_NEXTPTR   	32'h0131	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF3_AER_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF3_ARI_CAP_NEXTPTR   	32'h0132	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF3_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF3_ARI_CAP_NEXT_FUNC   	32'h0133	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_ARI_CAP_NEXT_FUNC_SZ	8

`define PCIE40E4__PF3_BAR0_APERTURE_SIZE   	32'h0134	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_BAR0_CONTROL   	32'h0135	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF3_BAR1_APERTURE_SIZE   	32'h0136	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_BAR1_CONTROL   	32'h0137	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF3_BAR2_APERTURE_SIZE   	32'h0138	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_BAR2_CONTROL   	32'h0139	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF3_BAR3_APERTURE_SIZE   	32'h013a	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_BAR3_CONTROL   	32'h013b	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF3_BAR4_APERTURE_SIZE   	32'h013c	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_BAR4_CONTROL   	32'h013d	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF3_BAR5_APERTURE_SIZE   	32'h013e	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_BAR5_CONTROL   	32'h013f	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF3_CAPABILITY_POINTER   	32'h0140	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_CAPABILITY_POINTER_SZ	8

`define PCIE40E4__PF3_CLASS_CODE   	32'h0141	// Type=HEX; Min=24'h000000, Max=24'hffffff
`define PCIE40E4__PF3_CLASS_CODE_SZ	24

`define PCIE40E4__PF3_DEV_CAP_MAX_PAYLOAD_SIZE   	32'h0142	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_DEV_CAP_MAX_PAYLOAD_SIZE_SZ	3

`define PCIE40E4__PF3_DSN_CAP_NEXTPTR   	32'h0143	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF3_DSN_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF3_EXPANSION_ROM_APERTURE_SIZE   	32'h0144	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_EXPANSION_ROM_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_EXPANSION_ROM_ENABLE   	32'h0145	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF3_EXPANSION_ROM_ENABLE_SZ	40

`define PCIE40E4__PF3_INTERRUPT_PIN   	32'h0146	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_INTERRUPT_PIN_SZ	3

`define PCIE40E4__PF3_MSIX_CAP_NEXTPTR   	32'h0147	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF3_MSIX_CAP_PBA_BIR   	32'h0148	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF3_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__PF3_MSIX_CAP_PBA_OFFSET   	32'h0149	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF3_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__PF3_MSIX_CAP_TABLE_BIR   	32'h014a	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF3_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__PF3_MSIX_CAP_TABLE_OFFSET   	32'h014b	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__PF3_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__PF3_MSIX_CAP_TABLE_SIZE   	32'h014c	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__PF3_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__PF3_MSI_CAP_MULTIMSGCAP   	32'h014d	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__PF3_MSI_CAP_MULTIMSGCAP_SZ	32

`define PCIE40E4__PF3_MSI_CAP_NEXTPTR   	32'h014e	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_MSI_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF3_MSI_CAP_PERVECMASKCAP   	32'h014f	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF3_MSI_CAP_PERVECMASKCAP_SZ	40

`define PCIE40E4__PF3_PCIE_CAP_NEXTPTR   	32'h0150	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF3_PM_CAP_NEXTPTR   	32'h0151	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PF3_PM_CAP_NEXTPTR_SZ	8

`define PCIE40E4__PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED   	32'h0152	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ	40

`define PCIE40E4__PF3_SRIOV_BAR0_APERTURE_SIZE   	32'h0153	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_SRIOV_BAR0_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_SRIOV_BAR0_CONTROL   	32'h0154	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR0_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_BAR1_APERTURE_SIZE   	32'h0155	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_SRIOV_BAR1_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_SRIOV_BAR1_CONTROL   	32'h0156	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR1_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_BAR2_APERTURE_SIZE   	32'h0157	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_SRIOV_BAR2_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_SRIOV_BAR2_CONTROL   	32'h0158	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR2_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_BAR3_APERTURE_SIZE   	32'h0159	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_SRIOV_BAR3_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_SRIOV_BAR3_CONTROL   	32'h015a	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR3_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_BAR4_APERTURE_SIZE   	32'h015b	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PF3_SRIOV_BAR4_APERTURE_SIZE_SZ	6

`define PCIE40E4__PF3_SRIOV_BAR4_CONTROL   	32'h015c	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR4_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_BAR5_APERTURE_SIZE   	32'h015d	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PF3_SRIOV_BAR5_APERTURE_SIZE_SZ	5

`define PCIE40E4__PF3_SRIOV_BAR5_CONTROL   	32'h015e	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_SRIOV_BAR5_CONTROL_SZ	3

`define PCIE40E4__PF3_SRIOV_CAP_INITIAL_VF   	32'h015f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF3_SRIOV_CAP_INITIAL_VF_SZ	16

`define PCIE40E4__PF3_SRIOV_CAP_NEXTPTR   	32'h0160	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF3_SRIOV_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF3_SRIOV_CAP_TOTAL_VF   	32'h0161	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF3_SRIOV_CAP_TOTAL_VF_SZ	16

`define PCIE40E4__PF3_SRIOV_CAP_VER   	32'h0162	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PF3_SRIOV_CAP_VER_SZ	4

`define PCIE40E4__PF3_SRIOV_FIRST_VF_OFFSET   	32'h0163	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF3_SRIOV_FIRST_VF_OFFSET_SZ	16

`define PCIE40E4__PF3_SRIOV_FUNC_DEP_LINK   	32'h0164	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF3_SRIOV_FUNC_DEP_LINK_SZ	16

`define PCIE40E4__PF3_SRIOV_SUPPORTED_PAGE_SIZE   	32'h0165	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PF3_SRIOV_SUPPORTED_PAGE_SIZE_SZ	32

`define PCIE40E4__PF3_SRIOV_VF_DEVICE_ID   	32'h0166	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PF3_SRIOV_VF_DEVICE_ID_SZ	16

`define PCIE40E4__PF3_TPHR_CAP_NEXTPTR   	32'h0167	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__PF3_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__PF3_TPHR_CAP_ST_MODE_SEL   	32'h0168	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__PF3_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__PL_CFG_STATE_ROBUSTNESS_ENABLE   	32'h0169	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_CFG_STATE_ROBUSTNESS_ENABLE_SZ	40

`define PCIE40E4__PL_DEEMPH_SOURCE_SELECT   	32'h016a	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_DEEMPH_SOURCE_SELECT_SZ	40

`define PCIE40E4__PL_DESKEW_ON_SKIP_IN_GEN12   	32'h016b	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DESKEW_ON_SKIP_IN_GEN12_SZ	40

`define PCIE40E4__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3   	32'h016c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_SZ	40

`define PCIE40E4__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4   	32'h016d	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4_SZ	40

`define PCIE40E4__PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2   	32'h016e	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_SZ	40

`define PCIE40E4__PL_DISABLE_DC_BALANCE   	32'h016f	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_DC_BALANCE_SZ	40

`define PCIE40E4__PL_DISABLE_EI_INFER_IN_L0   	32'h0170	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_EI_INFER_IN_L0_SZ	40

`define PCIE40E4__PL_DISABLE_LANE_REVERSAL   	32'h0171	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_LANE_REVERSAL_SZ	40

`define PCIE40E4__PL_DISABLE_LFSR_UPDATE_ON_SKP   	32'h0172	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_DISABLE_LFSR_UPDATE_ON_SKP_SZ	2

`define PCIE40E4__PL_DISABLE_RETRAIN_ON_EB_ERROR   	32'h0173	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_RETRAIN_ON_EB_ERROR_SZ	40

`define PCIE40E4__PL_DISABLE_RETRAIN_ON_FRAMING_ERROR   	32'h0174	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_SZ	40

`define PCIE40E4__PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR   	32'h0175	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR_SZ	16

`define PCIE40E4__PL_DISABLE_UPCONFIG_CAPABLE   	32'h0176	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_DISABLE_UPCONFIG_CAPABLE_SZ	40

`define PCIE40E4__PL_EQ_ADAPT_DISABLE_COEFF_CHECK   	32'h0177	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_ADAPT_DISABLE_COEFF_CHECK_SZ	2

`define PCIE40E4__PL_EQ_ADAPT_DISABLE_PRESET_CHECK   	32'h0178	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_ADAPT_DISABLE_PRESET_CHECK_SZ	2

`define PCIE40E4__PL_EQ_ADAPT_ITER_COUNT   	32'h0179	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PL_EQ_ADAPT_ITER_COUNT_SZ	5

`define PCIE40E4__PL_EQ_ADAPT_REJECT_RETRY_COUNT   	32'h017a	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_ADAPT_REJECT_RETRY_COUNT_SZ	2

`define PCIE40E4__PL_EQ_BYPASS_PHASE23   	32'h017b	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_BYPASS_PHASE23_SZ	2

`define PCIE40E4__PL_EQ_DEFAULT_RX_PRESET_HINT   	32'h017c	// Type=HEX; Min=6'h00, Max=6'h3f
`define PCIE40E4__PL_EQ_DEFAULT_RX_PRESET_HINT_SZ	6

`define PCIE40E4__PL_EQ_DEFAULT_TX_PRESET   	32'h017d	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PL_EQ_DEFAULT_TX_PRESET_SZ	8

`define PCIE40E4__PL_EQ_DISABLE_MISMATCH_CHECK   	32'h017e	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_EQ_DISABLE_MISMATCH_CHECK_SZ	40

`define PCIE40E4__PL_EQ_RX_ADAPT_EQ_PHASE0   	32'h017f	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_RX_ADAPT_EQ_PHASE0_SZ	2

`define PCIE40E4__PL_EQ_RX_ADAPT_EQ_PHASE1   	32'h0180	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_EQ_RX_ADAPT_EQ_PHASE1_SZ	2

`define PCIE40E4__PL_EQ_SHORT_ADAPT_PHASE   	32'h0181	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_EQ_SHORT_ADAPT_PHASE_SZ	40

`define PCIE40E4__PL_EQ_TX_8G_EQ_TS2_ENABLE   	32'h0182	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_EQ_TX_8G_EQ_TS2_ENABLE_SZ	40

`define PCIE40E4__PL_EXIT_LOOPBACK_ON_EI_ENTRY   	32'h0183	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_EXIT_LOOPBACK_ON_EI_ENTRY_SZ	40

`define PCIE40E4__PL_INFER_EI_DISABLE_LPBK_ACTIVE   	32'h0184	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_INFER_EI_DISABLE_LPBK_ACTIVE_SZ	40

`define PCIE40E4__PL_INFER_EI_DISABLE_REC_RC   	32'h0185	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_INFER_EI_DISABLE_REC_RC_SZ	40

`define PCIE40E4__PL_INFER_EI_DISABLE_REC_SPD   	32'h0186	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_INFER_EI_DISABLE_REC_SPD_SZ	40

`define PCIE40E4__PL_LANE0_EQ_CONTROL   	32'h0187	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE0_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE10_EQ_CONTROL   	32'h0188	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE10_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE11_EQ_CONTROL   	32'h0189	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE11_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE12_EQ_CONTROL   	32'h018a	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE12_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE13_EQ_CONTROL   	32'h018b	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE13_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE14_EQ_CONTROL   	32'h018c	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE14_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE15_EQ_CONTROL   	32'h018d	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE15_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE1_EQ_CONTROL   	32'h018e	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE1_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE2_EQ_CONTROL   	32'h018f	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE2_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE3_EQ_CONTROL   	32'h0190	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE3_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE4_EQ_CONTROL   	32'h0191	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE4_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE5_EQ_CONTROL   	32'h0192	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE5_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE6_EQ_CONTROL   	32'h0193	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE6_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE7_EQ_CONTROL   	32'h0194	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE7_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE8_EQ_CONTROL   	32'h0195	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE8_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LANE9_EQ_CONTROL   	32'h0196	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PL_LANE9_EQ_CONTROL_SZ	32

`define PCIE40E4__PL_LINK_CAP_MAX_LINK_SPEED   	32'h0197	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PL_LINK_CAP_MAX_LINK_SPEED_SZ	4

`define PCIE40E4__PL_LINK_CAP_MAX_LINK_WIDTH   	32'h0198	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__PL_LINK_CAP_MAX_LINK_WIDTH_SZ	5

`define PCIE40E4__PL_N_FTS   	32'h0199	// Type=DECIMAL; Min=0, Max=255
`define PCIE40E4__PL_N_FTS_SZ	32

`define PCIE40E4__PL_QUIESCE_GUARANTEE_DISABLE   	32'h019a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_QUIESCE_GUARANTEE_DISABLE_SZ	40

`define PCIE40E4__PL_REDO_EQ_SOURCE_SELECT   	32'h019b	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_REDO_EQ_SOURCE_SELECT_SZ	40

`define PCIE40E4__PL_REPORT_ALL_PHY_ERRORS   	32'h019c	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__PL_REPORT_ALL_PHY_ERRORS_SZ	8

`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS   	32'h019d	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS_SZ	2

`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_GEN3   	32'h019e	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_GEN3_SZ	4

`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_GEN4   	32'h019f	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PL_RX_ADAPT_TIMER_CLWS_GEN4_SZ	4

`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS   	32'h01a0	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS_SZ	2

`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_GEN3   	32'h01a1	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_GEN3_SZ	4

`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_GEN4   	32'h01a2	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__PL_RX_ADAPT_TIMER_RRL_GEN4_SZ	4

`define PCIE40E4__PL_RX_L0S_EXIT_TO_RECOVERY   	32'h01a3	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_RX_L0S_EXIT_TO_RECOVERY_SZ	2

`define PCIE40E4__PL_SIM_FAST_LINK_TRAINING   	32'h01a4	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__PL_SIM_FAST_LINK_TRAINING_SZ	2

`define PCIE40E4__PL_SRIS_ENABLE   	32'h01a5	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PL_SRIS_ENABLE_SZ	40

`define PCIE40E4__PL_SRIS_SKPOS_GEN_SPD_VEC   	32'h01a6	// Type=HEX; Min=7'h00, Max=7'h7f
`define PCIE40E4__PL_SRIS_SKPOS_GEN_SPD_VEC_SZ	7

`define PCIE40E4__PL_SRIS_SKPOS_REC_SPD_VEC   	32'h01a7	// Type=HEX; Min=7'h00, Max=7'h7f
`define PCIE40E4__PL_SRIS_SKPOS_REC_SPD_VEC_SZ	7

`define PCIE40E4__PL_UPSTREAM_FACING   	32'h01a8	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PL_UPSTREAM_FACING_SZ	40

`define PCIE40E4__PL_USER_SPARE   	32'h01a9	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PL_USER_SPARE_SZ	16

`define PCIE40E4__PM_ASPML0S_TIMEOUT   	32'h01aa	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PM_ASPML0S_TIMEOUT_SZ	16

`define PCIE40E4__PM_ASPML1_ENTRY_DELAY   	32'h01ab	// Type=HEX; Min=20'h00000, Max=20'hfffff
`define PCIE40E4__PM_ASPML1_ENTRY_DELAY_SZ	20

`define PCIE40E4__PM_ENABLE_L23_ENTRY   	32'h01ac	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__PM_ENABLE_L23_ENTRY_SZ	40

`define PCIE40E4__PM_ENABLE_SLOT_POWER_CAPTURE   	32'h01ad	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__PM_ENABLE_SLOT_POWER_CAPTURE_SZ	40

`define PCIE40E4__PM_L1_REENTRY_DELAY   	32'h01ae	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__PM_L1_REENTRY_DELAY_SZ	32

`define PCIE40E4__PM_PME_SERVICE_TIMEOUT_DELAY   	32'h01af	// Type=HEX; Min=20'h00000, Max=20'hfffff
`define PCIE40E4__PM_PME_SERVICE_TIMEOUT_DELAY_SZ	20

`define PCIE40E4__PM_PME_TURNOFF_ACK_DELAY   	32'h01b0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__PM_PME_TURNOFF_ACK_DELAY_SZ	16

`define PCIE40E4__SIM_DEVICE   	32'h01b1	// Type=STRING; Values=ULTRASCALE_PLUS,ULTRASCALE_PLUS_ES1,ULTRASCALE_PLUS_ES2
`define PCIE40E4__SIM_DEVICE_SZ	152

`define PCIE40E4__SIM_JTAG_IDCODE   	32'h01b2	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__SIM_JTAG_IDCODE_SZ	32

`define PCIE40E4__SIM_VERSION   	32'h01b3	// Type=STRING; Values=1.0,1.1,1.2,1.3,2.0,3.0,4.0
`define PCIE40E4__SIM_VERSION_SZ	24

`define PCIE40E4__SPARE_BIT0   	32'h01b4	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__SPARE_BIT0_SZ	40

`define PCIE40E4__SPARE_BIT1   	32'h01b5	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT1_SZ	32

`define PCIE40E4__SPARE_BIT2   	32'h01b6	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT2_SZ	32

`define PCIE40E4__SPARE_BIT3   	32'h01b7	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__SPARE_BIT3_SZ	40

`define PCIE40E4__SPARE_BIT4   	32'h01b8	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT4_SZ	32

`define PCIE40E4__SPARE_BIT5   	32'h01b9	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT5_SZ	32

`define PCIE40E4__SPARE_BIT6   	32'h01ba	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT6_SZ	32

`define PCIE40E4__SPARE_BIT7   	32'h01bb	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT7_SZ	32

`define PCIE40E4__SPARE_BIT8   	32'h01bc	// Type=DECIMAL; Values=0,1
`define PCIE40E4__SPARE_BIT8_SZ	32

`define PCIE40E4__SPARE_BYTE0   	32'h01bd	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__SPARE_BYTE0_SZ	8

`define PCIE40E4__SPARE_BYTE1   	32'h01be	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__SPARE_BYTE1_SZ	8

`define PCIE40E4__SPARE_BYTE2   	32'h01bf	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__SPARE_BYTE2_SZ	8

`define PCIE40E4__SPARE_BYTE3   	32'h01c0	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__SPARE_BYTE3_SZ	8

`define PCIE40E4__SPARE_WORD0   	32'h01c1	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__SPARE_WORD0_SZ	32

`define PCIE40E4__SPARE_WORD1   	32'h01c2	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__SPARE_WORD1_SZ	32

`define PCIE40E4__SPARE_WORD2   	32'h01c3	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__SPARE_WORD2_SZ	32

`define PCIE40E4__SPARE_WORD3   	32'h01c4	// Type=HEX; Min=32'h00000000, Max=32'hffffffff
`define PCIE40E4__SPARE_WORD3_SZ	32

`define PCIE40E4__SRIOV_CAP_ENABLE   	32'h01c5	// Type=HEX; Min=4'h0, Max=4'hf
`define PCIE40E4__SRIOV_CAP_ENABLE_SZ	4

`define PCIE40E4__TL2CFG_IF_PARITY_CHK   	32'h01c6	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__TL2CFG_IF_PARITY_CHK_SZ	40

`define PCIE40E4__TL_COMPLETION_RAM_NUM_TLPS   	32'h01c7	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__TL_COMPLETION_RAM_NUM_TLPS_SZ	2

`define PCIE40E4__TL_COMPLETION_RAM_SIZE   	32'h01c8	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__TL_COMPLETION_RAM_SIZE_SZ	2

`define PCIE40E4__TL_CREDITS_CD   	32'h01c9	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__TL_CREDITS_CD_SZ	12

`define PCIE40E4__TL_CREDITS_CH   	32'h01ca	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__TL_CREDITS_CH_SZ	8

`define PCIE40E4__TL_CREDITS_NPD   	32'h01cb	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__TL_CREDITS_NPD_SZ	12

`define PCIE40E4__TL_CREDITS_NPH   	32'h01cc	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__TL_CREDITS_NPH_SZ	8

`define PCIE40E4__TL_CREDITS_PD   	32'h01cd	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__TL_CREDITS_PD_SZ	12

`define PCIE40E4__TL_CREDITS_PH   	32'h01ce	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__TL_CREDITS_PH_SZ	8

`define PCIE40E4__TL_FC_UPDATE_MIN_INTERVAL_TIME   	32'h01cf	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__TL_FC_UPDATE_MIN_INTERVAL_TIME_SZ	5

`define PCIE40E4__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT   	32'h01d0	// Type=HEX; Min=5'h00, Max=5'h1f
`define PCIE40E4__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT_SZ	5

`define PCIE40E4__TL_PF_ENABLE_REG   	32'h01d1	// Type=HEX; Min=2'h0, Max=2'h3
`define PCIE40E4__TL_PF_ENABLE_REG_SZ	2

`define PCIE40E4__TL_POSTED_RAM_SIZE   	32'h01d2	// Type=HEX; Min=1'h0, Max=1'h1
`define PCIE40E4__TL_POSTED_RAM_SIZE_SZ	1

`define PCIE40E4__TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE   	32'h01d3	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE_SZ	40

`define PCIE40E4__TL_RX_COMPLETION_TO_RAM_READ_PIPELINE   	32'h01d4	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_COMPLETION_TO_RAM_READ_PIPELINE_SZ	40

`define PCIE40E4__TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE   	32'h01d5	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE_SZ	40

`define PCIE40E4__TL_RX_POSTED_FROM_RAM_READ_PIPELINE   	32'h01d6	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_POSTED_FROM_RAM_READ_PIPELINE_SZ	40

`define PCIE40E4__TL_RX_POSTED_TO_RAM_READ_PIPELINE   	32'h01d7	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_POSTED_TO_RAM_READ_PIPELINE_SZ	40

`define PCIE40E4__TL_RX_POSTED_TO_RAM_WRITE_PIPELINE   	32'h01d8	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_RX_POSTED_TO_RAM_WRITE_PIPELINE_SZ	40

`define PCIE40E4__TL_TX_MUX_STRICT_PRIORITY   	32'h01d9	// Type=BOOLSTRING; Values=TRUE,FALSE
`define PCIE40E4__TL_TX_MUX_STRICT_PRIORITY_SZ	40

`define PCIE40E4__TL_TX_TLP_STRADDLE_ENABLE   	32'h01da	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_TX_TLP_STRADDLE_ENABLE_SZ	40

`define PCIE40E4__TL_TX_TLP_TERMINATE_PARITY   	32'h01db	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TL_TX_TLP_TERMINATE_PARITY_SZ	40

`define PCIE40E4__TL_USER_SPARE   	32'h01dc	// Type=HEX; Min=16'h0000, Max=16'hffff
`define PCIE40E4__TL_USER_SPARE_SZ	16

`define PCIE40E4__TPH_FROM_RAM_PIPELINE   	32'h01dd	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TPH_FROM_RAM_PIPELINE_SZ	40

`define PCIE40E4__TPH_TO_RAM_PIPELINE   	32'h01de	// Type=BOOLSTRING; Values=FALSE,TRUE
`define PCIE40E4__TPH_TO_RAM_PIPELINE_SZ	40

`define PCIE40E4__VF0_CAPABILITY_POINTER   	32'h01df	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VF0_CAPABILITY_POINTER_SZ	8

`define PCIE40E4__VFG0_ARI_CAP_NEXTPTR   	32'h01e0	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG0_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG0_MSIX_CAP_NEXTPTR   	32'h01e1	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG0_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG0_MSIX_CAP_PBA_BIR   	32'h01e2	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG0_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__VFG0_MSIX_CAP_PBA_OFFSET   	32'h01e3	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG0_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__VFG0_MSIX_CAP_TABLE_BIR   	32'h01e4	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG0_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__VFG0_MSIX_CAP_TABLE_OFFSET   	32'h01e5	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG0_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__VFG0_MSIX_CAP_TABLE_SIZE   	32'h01e6	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__VFG0_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__VFG0_PCIE_CAP_NEXTPTR   	32'h01e7	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG0_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG0_TPHR_CAP_NEXTPTR   	32'h01e8	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG0_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG0_TPHR_CAP_ST_MODE_SEL   	32'h01e9	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__VFG0_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__VFG1_ARI_CAP_NEXTPTR   	32'h01ea	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG1_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG1_MSIX_CAP_NEXTPTR   	32'h01eb	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG1_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG1_MSIX_CAP_PBA_BIR   	32'h01ec	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG1_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__VFG1_MSIX_CAP_PBA_OFFSET   	32'h01ed	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG1_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__VFG1_MSIX_CAP_TABLE_BIR   	32'h01ee	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG1_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__VFG1_MSIX_CAP_TABLE_OFFSET   	32'h01ef	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG1_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__VFG1_MSIX_CAP_TABLE_SIZE   	32'h01f0	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__VFG1_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__VFG1_PCIE_CAP_NEXTPTR   	32'h01f1	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG1_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG1_TPHR_CAP_NEXTPTR   	32'h01f2	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG1_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG1_TPHR_CAP_ST_MODE_SEL   	32'h01f3	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__VFG1_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__VFG2_ARI_CAP_NEXTPTR   	32'h01f4	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG2_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG2_MSIX_CAP_NEXTPTR   	32'h01f5	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG2_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG2_MSIX_CAP_PBA_BIR   	32'h01f6	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG2_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__VFG2_MSIX_CAP_PBA_OFFSET   	32'h01f7	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG2_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__VFG2_MSIX_CAP_TABLE_BIR   	32'h01f8	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG2_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__VFG2_MSIX_CAP_TABLE_OFFSET   	32'h01f9	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG2_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__VFG2_MSIX_CAP_TABLE_SIZE   	32'h01fa	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__VFG2_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__VFG2_PCIE_CAP_NEXTPTR   	32'h01fb	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG2_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG2_TPHR_CAP_NEXTPTR   	32'h01fc	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG2_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG2_TPHR_CAP_ST_MODE_SEL   	32'h01fd	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__VFG2_TPHR_CAP_ST_MODE_SEL_SZ	3

`define PCIE40E4__VFG3_ARI_CAP_NEXTPTR   	32'h01fe	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG3_ARI_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG3_MSIX_CAP_NEXTPTR   	32'h01ff	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG3_MSIX_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG3_MSIX_CAP_PBA_BIR   	32'h0200	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG3_MSIX_CAP_PBA_BIR_SZ	32

`define PCIE40E4__VFG3_MSIX_CAP_PBA_OFFSET   	32'h0201	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG3_MSIX_CAP_PBA_OFFSET_SZ	29

`define PCIE40E4__VFG3_MSIX_CAP_TABLE_BIR   	32'h0202	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7
`define PCIE40E4__VFG3_MSIX_CAP_TABLE_BIR_SZ	32

`define PCIE40E4__VFG3_MSIX_CAP_TABLE_OFFSET   	32'h0203	// Type=HEX; Min=29'h00000000, Max=29'h1fffffff
`define PCIE40E4__VFG3_MSIX_CAP_TABLE_OFFSET_SZ	29

`define PCIE40E4__VFG3_MSIX_CAP_TABLE_SIZE   	32'h0204	// Type=HEX; Min=11'h000, Max=11'h7ff
`define PCIE40E4__VFG3_MSIX_CAP_TABLE_SIZE_SZ	11

`define PCIE40E4__VFG3_PCIE_CAP_NEXTPTR   	32'h0205	// Type=HEX; Min=8'h00, Max=8'hff
`define PCIE40E4__VFG3_PCIE_CAP_NEXTPTR_SZ	8

`define PCIE40E4__VFG3_TPHR_CAP_NEXTPTR   	32'h0206	// Type=HEX; Min=12'h000, Max=12'hfff
`define PCIE40E4__VFG3_TPHR_CAP_NEXTPTR_SZ	12

`define PCIE40E4__VFG3_TPHR_CAP_ST_MODE_SEL   	32'h0207	// Type=HEX; Min=3'h0, Max=3'h7
`define PCIE40E4__VFG3_TPHR_CAP_ST_MODE_SEL_SZ	3

`endif  // B_PCIE40E4_DEFINES_VH
