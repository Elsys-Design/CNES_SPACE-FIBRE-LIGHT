// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_FP_SRCMX_OPTINV_DEFINES_VH
`else
`define B_DSP_FP_SRCMX_OPTINV_DEFINES_VH

// Look-up table parameters
//

`define DSP_FP_SRCMX_OPTINV_ADDR_N  3
`define DSP_FP_SRCMX_OPTINV_ADDR_SZ 32
`define DSP_FP_SRCMX_OPTINV_DATA_SZ 1

// Attribute addresses
//

`define DSP_FP_SRCMX_OPTINV__IS_ASYNC_RST_INVERTED    32'h00000000
`define DSP_FP_SRCMX_OPTINV__IS_ASYNC_RST_INVERTED_SZ 1

`define DSP_FP_SRCMX_OPTINV__IS_CLK_INVERTED    32'h00000001
`define DSP_FP_SRCMX_OPTINV__IS_CLK_INVERTED_SZ 1

`define DSP_FP_SRCMX_OPTINV__IS_RSTD_INVERTED    32'h00000002
`define DSP_FP_SRCMX_OPTINV__IS_RSTD_INVERTED_SZ 1

`endif  // B_DSP_FP_SRCMX_OPTINV_DEFINES_VH