// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTME5_QUAD_DEFINES_VH
`else
`define B_GTME5_QUAD_DEFINES_VH

// Look-up table parameters
//

`define GTME5_QUAD_ADDR_N  648
`define GTME5_QUAD_ADDR_SZ 32
`define GTME5_QUAD_DATA_SZ 192

// Attribute addresses
//

`define GTME5_QUAD__A_CFG0    32'h00000000
`define GTME5_QUAD__A_CFG0_SZ 32

`define GTME5_QUAD__A_CFG1    32'h00000001
`define GTME5_QUAD__A_CFG1_SZ 32

`define GTME5_QUAD__A_CFG2    32'h00000002
`define GTME5_QUAD__A_CFG2_SZ 32

`define GTME5_QUAD__A_CFG3    32'h00000003
`define GTME5_QUAD__A_CFG3_SZ 32

`define GTME5_QUAD__A_CFG4    32'h00000004
`define GTME5_QUAD__A_CFG4_SZ 32

`define GTME5_QUAD__A_CFG5    32'h00000005
`define GTME5_QUAD__A_CFG5_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG0    32'h00000006
`define GTME5_QUAD__CH0_CHCLK_CFG0_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG1    32'h00000007
`define GTME5_QUAD__CH0_CHCLK_CFG1_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG2    32'h00000008
`define GTME5_QUAD__CH0_CHCLK_CFG2_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG3    32'h00000009
`define GTME5_QUAD__CH0_CHCLK_CFG3_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG4    32'h0000000a
`define GTME5_QUAD__CH0_CHCLK_CFG4_SZ 32

`define GTME5_QUAD__CH0_CHCLK_CFG5    32'h0000000b
`define GTME5_QUAD__CH0_CHCLK_CFG5_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG0    32'h0000000c
`define GTME5_QUAD__CH0_EYESCAN_CFG0_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG1    32'h0000000d
`define GTME5_QUAD__CH0_EYESCAN_CFG1_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG2    32'h0000000e
`define GTME5_QUAD__CH0_EYESCAN_CFG2_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG3    32'h0000000f
`define GTME5_QUAD__CH0_EYESCAN_CFG3_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG4    32'h00000010
`define GTME5_QUAD__CH0_EYESCAN_CFG4_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG5    32'h00000011
`define GTME5_QUAD__CH0_EYESCAN_CFG5_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG6    32'h00000012
`define GTME5_QUAD__CH0_EYESCAN_CFG6_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG7    32'h00000013
`define GTME5_QUAD__CH0_EYESCAN_CFG7_SZ 32

`define GTME5_QUAD__CH0_EYESCAN_CFG8    32'h00000014
`define GTME5_QUAD__CH0_EYESCAN_CFG8_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG0    32'h00000015
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG0_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG1    32'h00000016
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG1_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG2    32'h00000017
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG2_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG3    32'h00000018
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG3_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG4    32'h00000019
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG4_SZ 32

`define GTME5_QUAD__CH0_FABRIC_INTF_CFG5    32'h0000001a
`define GTME5_QUAD__CH0_FABRIC_INTF_CFG5_SZ 32

`define GTME5_QUAD__CH0_INSTANTIATED    32'h0000001b
`define GTME5_QUAD__CH0_INSTANTIATED_SZ 1

`define GTME5_QUAD__CH0_MONITOR_CFG0    32'h0000001c
`define GTME5_QUAD__CH0_MONITOR_CFG0_SZ 32

`define GTME5_QUAD__CH0_PMA_MISC_CFG0    32'h0000001d
`define GTME5_QUAD__CH0_PMA_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH0_RESET_BYP_HDSHK_CFG    32'h0000001e
`define GTME5_QUAD__CH0_RESET_BYP_HDSHK_CFG_SZ 32

`define GTME5_QUAD__CH0_RESET_CFG    32'h0000001f
`define GTME5_QUAD__CH0_RESET_CFG_SZ 32

`define GTME5_QUAD__CH0_RESET_LOOPER_ID_CFG    32'h00000020
`define GTME5_QUAD__CH0_RESET_LOOPER_ID_CFG_SZ 32

`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG0    32'h00000021
`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG0_SZ 32

`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG1    32'h00000022
`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG1_SZ 32

`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG2    32'h00000023
`define GTME5_QUAD__CH0_RESET_LOOP_ID_CFG2_SZ 32

`define GTME5_QUAD__CH0_RESET_TIME_CFG0    32'h00000024
`define GTME5_QUAD__CH0_RESET_TIME_CFG0_SZ 32

`define GTME5_QUAD__CH0_RESET_TIME_CFG1    32'h00000025
`define GTME5_QUAD__CH0_RESET_TIME_CFG1_SZ 32

`define GTME5_QUAD__CH0_RESET_TIME_CFG2    32'h00000026
`define GTME5_QUAD__CH0_RESET_TIME_CFG2_SZ 32

`define GTME5_QUAD__CH0_RESET_TIME_CFG3    32'h00000027
`define GTME5_QUAD__CH0_RESET_TIME_CFG3_SZ 32

`define GTME5_QUAD__CH0_RXOUTCLK_FREQ    32'h00000028
`define GTME5_QUAD__CH0_RXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH0_RXOUTCLK_REF_FREQ    32'h00000029
`define GTME5_QUAD__CH0_RXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH0_RXOUTCLK_REF_SOURCE    32'h0000002a
`define GTME5_QUAD__CH0_RXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH0_RX_APT_CFG0    32'h0000002b
`define GTME5_QUAD__CH0_RX_APT_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG1    32'h0000002c
`define GTME5_QUAD__CH0_RX_APT_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG10    32'h0000002d
`define GTME5_QUAD__CH0_RX_APT_CFG10_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG11    32'h0000002e
`define GTME5_QUAD__CH0_RX_APT_CFG11_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG12    32'h0000002f
`define GTME5_QUAD__CH0_RX_APT_CFG12_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG13    32'h00000030
`define GTME5_QUAD__CH0_RX_APT_CFG13_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG14    32'h00000031
`define GTME5_QUAD__CH0_RX_APT_CFG14_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG15    32'h00000032
`define GTME5_QUAD__CH0_RX_APT_CFG15_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG16    32'h00000033
`define GTME5_QUAD__CH0_RX_APT_CFG16_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG17    32'h00000034
`define GTME5_QUAD__CH0_RX_APT_CFG17_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG18    32'h00000035
`define GTME5_QUAD__CH0_RX_APT_CFG18_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG19    32'h00000036
`define GTME5_QUAD__CH0_RX_APT_CFG19_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG2    32'h00000037
`define GTME5_QUAD__CH0_RX_APT_CFG2_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG20    32'h00000038
`define GTME5_QUAD__CH0_RX_APT_CFG20_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG21    32'h00000039
`define GTME5_QUAD__CH0_RX_APT_CFG21_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG22    32'h0000003a
`define GTME5_QUAD__CH0_RX_APT_CFG22_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG23    32'h0000003b
`define GTME5_QUAD__CH0_RX_APT_CFG23_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG24    32'h0000003c
`define GTME5_QUAD__CH0_RX_APT_CFG24_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG25    32'h0000003d
`define GTME5_QUAD__CH0_RX_APT_CFG25_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG26    32'h0000003e
`define GTME5_QUAD__CH0_RX_APT_CFG26_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG27    32'h0000003f
`define GTME5_QUAD__CH0_RX_APT_CFG27_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG28    32'h00000040
`define GTME5_QUAD__CH0_RX_APT_CFG28_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG29    32'h00000041
`define GTME5_QUAD__CH0_RX_APT_CFG29_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG3    32'h00000042
`define GTME5_QUAD__CH0_RX_APT_CFG3_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG30    32'h00000043
`define GTME5_QUAD__CH0_RX_APT_CFG30_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG31    32'h00000044
`define GTME5_QUAD__CH0_RX_APT_CFG31_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG32    32'h00000045
`define GTME5_QUAD__CH0_RX_APT_CFG32_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG33    32'h00000046
`define GTME5_QUAD__CH0_RX_APT_CFG33_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG34    32'h00000047
`define GTME5_QUAD__CH0_RX_APT_CFG34_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG35    32'h00000048
`define GTME5_QUAD__CH0_RX_APT_CFG35_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG36    32'h00000049
`define GTME5_QUAD__CH0_RX_APT_CFG36_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG37    32'h0000004a
`define GTME5_QUAD__CH0_RX_APT_CFG37_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG38    32'h0000004b
`define GTME5_QUAD__CH0_RX_APT_CFG38_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG39    32'h0000004c
`define GTME5_QUAD__CH0_RX_APT_CFG39_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG4    32'h0000004d
`define GTME5_QUAD__CH0_RX_APT_CFG4_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG40    32'h0000004e
`define GTME5_QUAD__CH0_RX_APT_CFG40_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG41    32'h0000004f
`define GTME5_QUAD__CH0_RX_APT_CFG41_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG42    32'h00000050
`define GTME5_QUAD__CH0_RX_APT_CFG42_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG43    32'h00000051
`define GTME5_QUAD__CH0_RX_APT_CFG43_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG44    32'h00000052
`define GTME5_QUAD__CH0_RX_APT_CFG44_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG45    32'h00000053
`define GTME5_QUAD__CH0_RX_APT_CFG45_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG46    32'h00000054
`define GTME5_QUAD__CH0_RX_APT_CFG46_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG47    32'h00000055
`define GTME5_QUAD__CH0_RX_APT_CFG47_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG48    32'h00000056
`define GTME5_QUAD__CH0_RX_APT_CFG48_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG49    32'h00000057
`define GTME5_QUAD__CH0_RX_APT_CFG49_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG5    32'h00000058
`define GTME5_QUAD__CH0_RX_APT_CFG5_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG50    32'h00000059
`define GTME5_QUAD__CH0_RX_APT_CFG50_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG51    32'h0000005a
`define GTME5_QUAD__CH0_RX_APT_CFG51_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG52    32'h0000005b
`define GTME5_QUAD__CH0_RX_APT_CFG52_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG53    32'h0000005c
`define GTME5_QUAD__CH0_RX_APT_CFG53_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG54    32'h0000005d
`define GTME5_QUAD__CH0_RX_APT_CFG54_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG55    32'h0000005e
`define GTME5_QUAD__CH0_RX_APT_CFG55_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG56    32'h0000005f
`define GTME5_QUAD__CH0_RX_APT_CFG56_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG57    32'h00000060
`define GTME5_QUAD__CH0_RX_APT_CFG57_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG58    32'h00000061
`define GTME5_QUAD__CH0_RX_APT_CFG58_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG6    32'h00000062
`define GTME5_QUAD__CH0_RX_APT_CFG6_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG7    32'h00000063
`define GTME5_QUAD__CH0_RX_APT_CFG7_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG8    32'h00000064
`define GTME5_QUAD__CH0_RX_APT_CFG8_SZ 32

`define GTME5_QUAD__CH0_RX_APT_CFG9    32'h00000065
`define GTME5_QUAD__CH0_RX_APT_CFG9_SZ 32

`define GTME5_QUAD__CH0_RX_CAL_CFG0    32'h00000066
`define GTME5_QUAD__CH0_RX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_CAL_CFG1    32'h00000067
`define GTME5_QUAD__CH0_RX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_CAL_CFG2    32'h00000068
`define GTME5_QUAD__CH0_RX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG0    32'h00000069
`define GTME5_QUAD__CH0_RX_CDR_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG1    32'h0000006a
`define GTME5_QUAD__CH0_RX_CDR_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG2    32'h0000006b
`define GTME5_QUAD__CH0_RX_CDR_CFG2_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG3    32'h0000006c
`define GTME5_QUAD__CH0_RX_CDR_CFG3_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG4    32'h0000006d
`define GTME5_QUAD__CH0_RX_CDR_CFG4_SZ 32

`define GTME5_QUAD__CH0_RX_CDR_CFG5    32'h0000006e
`define GTME5_QUAD__CH0_RX_CDR_CFG5_SZ 32

`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG0    32'h0000006f
`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG1    32'h00000070
`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG2    32'h00000071
`define GTME5_QUAD__CH0_RX_CTLE_ADC_CFG2_SZ 32

`define GTME5_QUAD__CH0_RX_CTLE_HF_CFG0    32'h00000072
`define GTME5_QUAD__CH0_RX_CTLE_HF_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_CTLE_HF_CFG1    32'h00000073
`define GTME5_QUAD__CH0_RX_CTLE_HF_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_DSP_CFG0    32'h00000074
`define GTME5_QUAD__CH0_RX_DSP_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_DSP_CFG1    32'h00000075
`define GTME5_QUAD__CH0_RX_DSP_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_MISC_CFG1    32'h00000076
`define GTME5_QUAD__CH0_RX_MISC_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_PAD_CFG0    32'h00000077
`define GTME5_QUAD__CH0_RX_PAD_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_PAD_CFG1    32'h00000078
`define GTME5_QUAD__CH0_RX_PAD_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_PCS_CFG0    32'h00000079
`define GTME5_QUAD__CH0_RX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_PCS_CFG1    32'h0000007a
`define GTME5_QUAD__CH0_RX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_RSV_CFG0    32'h0000007b
`define GTME5_QUAD__CH0_RX_RSV_CFG0_SZ 32

`define GTME5_QUAD__CH0_RX_RSV_CFG1    32'h0000007c
`define GTME5_QUAD__CH0_RX_RSV_CFG1_SZ 32

`define GTME5_QUAD__CH0_RX_SPARE_CFG0    32'h0000007d
`define GTME5_QUAD__CH0_RX_SPARE_CFG0_SZ 32

`define GTME5_QUAD__CH0_SIM_MODE    32'h0000007e
`define GTME5_QUAD__CH0_SIM_MODE_SZ 48

`define GTME5_QUAD__CH0_SIM_RECEIVER_DETECT_PASS    32'h0000007f
`define GTME5_QUAD__CH0_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTME5_QUAD__CH0_SIM_RESET_SPEEDUP    32'h00000080
`define GTME5_QUAD__CH0_SIM_RESET_SPEEDUP_SZ 40

`define GTME5_QUAD__CH0_TXOUTCLK_FREQ    32'h00000081
`define GTME5_QUAD__CH0_TXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH0_TXOUTCLK_REF_FREQ    32'h00000082
`define GTME5_QUAD__CH0_TXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH0_TXOUTCLK_REF_SOURCE    32'h00000083
`define GTME5_QUAD__CH0_TXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH0_TX_CAL_CFG0    32'h00000084
`define GTME5_QUAD__CH0_TX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH0_TX_CAL_CFG1    32'h00000085
`define GTME5_QUAD__CH0_TX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH0_TX_CAL_CFG2    32'h00000086
`define GTME5_QUAD__CH0_TX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH0_TX_CTRL_CFG0    32'h00000087
`define GTME5_QUAD__CH0_TX_CTRL_CFG0_SZ 32

`define GTME5_QUAD__CH0_TX_CTRL_CFG1    32'h00000088
`define GTME5_QUAD__CH0_TX_CTRL_CFG1_SZ 32

`define GTME5_QUAD__CH0_TX_CTRL_CFG2    32'h00000089
`define GTME5_QUAD__CH0_TX_CTRL_CFG2_SZ 32

`define GTME5_QUAD__CH0_TX_CTRL_CFG3    32'h0000008a
`define GTME5_QUAD__CH0_TX_CTRL_CFG3_SZ 32

`define GTME5_QUAD__CH0_TX_MISC_CFG0    32'h0000008b
`define GTME5_QUAD__CH0_TX_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG0    32'h0000008c
`define GTME5_QUAD__CH0_TX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG1    32'h0000008d
`define GTME5_QUAD__CH0_TX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG2    32'h0000008e
`define GTME5_QUAD__CH0_TX_PCS_CFG2_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG3    32'h0000008f
`define GTME5_QUAD__CH0_TX_PCS_CFG3_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG4    32'h00000090
`define GTME5_QUAD__CH0_TX_PCS_CFG4_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG5    32'h00000091
`define GTME5_QUAD__CH0_TX_PCS_CFG5_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG6    32'h00000092
`define GTME5_QUAD__CH0_TX_PCS_CFG6_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG7    32'h00000093
`define GTME5_QUAD__CH0_TX_PCS_CFG7_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG8    32'h00000094
`define GTME5_QUAD__CH0_TX_PCS_CFG8_SZ 32

`define GTME5_QUAD__CH0_TX_PCS_CFG9    32'h00000095
`define GTME5_QUAD__CH0_TX_PCS_CFG9_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG0    32'h00000096
`define GTME5_QUAD__CH1_CHCLK_CFG0_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG1    32'h00000097
`define GTME5_QUAD__CH1_CHCLK_CFG1_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG2    32'h00000098
`define GTME5_QUAD__CH1_CHCLK_CFG2_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG3    32'h00000099
`define GTME5_QUAD__CH1_CHCLK_CFG3_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG4    32'h0000009a
`define GTME5_QUAD__CH1_CHCLK_CFG4_SZ 32

`define GTME5_QUAD__CH1_CHCLK_CFG5    32'h0000009b
`define GTME5_QUAD__CH1_CHCLK_CFG5_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG0    32'h0000009c
`define GTME5_QUAD__CH1_EYESCAN_CFG0_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG1    32'h0000009d
`define GTME5_QUAD__CH1_EYESCAN_CFG1_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG2    32'h0000009e
`define GTME5_QUAD__CH1_EYESCAN_CFG2_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG3    32'h0000009f
`define GTME5_QUAD__CH1_EYESCAN_CFG3_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG4    32'h000000a0
`define GTME5_QUAD__CH1_EYESCAN_CFG4_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG5    32'h000000a1
`define GTME5_QUAD__CH1_EYESCAN_CFG5_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG6    32'h000000a2
`define GTME5_QUAD__CH1_EYESCAN_CFG6_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG7    32'h000000a3
`define GTME5_QUAD__CH1_EYESCAN_CFG7_SZ 32

`define GTME5_QUAD__CH1_EYESCAN_CFG8    32'h000000a4
`define GTME5_QUAD__CH1_EYESCAN_CFG8_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG0    32'h000000a5
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG0_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG1    32'h000000a6
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG1_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG2    32'h000000a7
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG2_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG3    32'h000000a8
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG3_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG4    32'h000000a9
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG4_SZ 32

`define GTME5_QUAD__CH1_FABRIC_INTF_CFG5    32'h000000aa
`define GTME5_QUAD__CH1_FABRIC_INTF_CFG5_SZ 32

`define GTME5_QUAD__CH1_INSTANTIATED    32'h000000ab
`define GTME5_QUAD__CH1_INSTANTIATED_SZ 1

`define GTME5_QUAD__CH1_MONITOR_CFG0    32'h000000ac
`define GTME5_QUAD__CH1_MONITOR_CFG0_SZ 32

`define GTME5_QUAD__CH1_PMA_MISC_CFG0    32'h000000ad
`define GTME5_QUAD__CH1_PMA_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH1_RESET_BYP_HDSHK_CFG    32'h000000ae
`define GTME5_QUAD__CH1_RESET_BYP_HDSHK_CFG_SZ 32

`define GTME5_QUAD__CH1_RESET_CFG    32'h000000af
`define GTME5_QUAD__CH1_RESET_CFG_SZ 32

`define GTME5_QUAD__CH1_RESET_LOOPER_ID_CFG    32'h000000b0
`define GTME5_QUAD__CH1_RESET_LOOPER_ID_CFG_SZ 32

`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG0    32'h000000b1
`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG0_SZ 32

`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG1    32'h000000b2
`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG1_SZ 32

`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG2    32'h000000b3
`define GTME5_QUAD__CH1_RESET_LOOP_ID_CFG2_SZ 32

`define GTME5_QUAD__CH1_RESET_TIME_CFG0    32'h000000b4
`define GTME5_QUAD__CH1_RESET_TIME_CFG0_SZ 32

`define GTME5_QUAD__CH1_RESET_TIME_CFG1    32'h000000b5
`define GTME5_QUAD__CH1_RESET_TIME_CFG1_SZ 32

`define GTME5_QUAD__CH1_RESET_TIME_CFG2    32'h000000b6
`define GTME5_QUAD__CH1_RESET_TIME_CFG2_SZ 32

`define GTME5_QUAD__CH1_RESET_TIME_CFG3    32'h000000b7
`define GTME5_QUAD__CH1_RESET_TIME_CFG3_SZ 32

`define GTME5_QUAD__CH1_RXOUTCLK_FREQ    32'h000000b8
`define GTME5_QUAD__CH1_RXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH1_RXOUTCLK_REF_FREQ    32'h000000b9
`define GTME5_QUAD__CH1_RXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH1_RXOUTCLK_REF_SOURCE    32'h000000ba
`define GTME5_QUAD__CH1_RXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH1_RX_APT_CFG0    32'h000000bb
`define GTME5_QUAD__CH1_RX_APT_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG1    32'h000000bc
`define GTME5_QUAD__CH1_RX_APT_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG10    32'h000000bd
`define GTME5_QUAD__CH1_RX_APT_CFG10_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG11    32'h000000be
`define GTME5_QUAD__CH1_RX_APT_CFG11_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG12    32'h000000bf
`define GTME5_QUAD__CH1_RX_APT_CFG12_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG13    32'h000000c0
`define GTME5_QUAD__CH1_RX_APT_CFG13_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG14    32'h000000c1
`define GTME5_QUAD__CH1_RX_APT_CFG14_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG15    32'h000000c2
`define GTME5_QUAD__CH1_RX_APT_CFG15_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG16    32'h000000c3
`define GTME5_QUAD__CH1_RX_APT_CFG16_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG17    32'h000000c4
`define GTME5_QUAD__CH1_RX_APT_CFG17_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG18    32'h000000c5
`define GTME5_QUAD__CH1_RX_APT_CFG18_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG19    32'h000000c6
`define GTME5_QUAD__CH1_RX_APT_CFG19_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG2    32'h000000c7
`define GTME5_QUAD__CH1_RX_APT_CFG2_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG20    32'h000000c8
`define GTME5_QUAD__CH1_RX_APT_CFG20_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG21    32'h000000c9
`define GTME5_QUAD__CH1_RX_APT_CFG21_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG22    32'h000000ca
`define GTME5_QUAD__CH1_RX_APT_CFG22_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG23    32'h000000cb
`define GTME5_QUAD__CH1_RX_APT_CFG23_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG24    32'h000000cc
`define GTME5_QUAD__CH1_RX_APT_CFG24_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG25    32'h000000cd
`define GTME5_QUAD__CH1_RX_APT_CFG25_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG26    32'h000000ce
`define GTME5_QUAD__CH1_RX_APT_CFG26_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG27    32'h000000cf
`define GTME5_QUAD__CH1_RX_APT_CFG27_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG28    32'h000000d0
`define GTME5_QUAD__CH1_RX_APT_CFG28_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG29    32'h000000d1
`define GTME5_QUAD__CH1_RX_APT_CFG29_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG3    32'h000000d2
`define GTME5_QUAD__CH1_RX_APT_CFG3_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG30    32'h000000d3
`define GTME5_QUAD__CH1_RX_APT_CFG30_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG31    32'h000000d4
`define GTME5_QUAD__CH1_RX_APT_CFG31_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG32    32'h000000d5
`define GTME5_QUAD__CH1_RX_APT_CFG32_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG33    32'h000000d6
`define GTME5_QUAD__CH1_RX_APT_CFG33_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG34    32'h000000d7
`define GTME5_QUAD__CH1_RX_APT_CFG34_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG35    32'h000000d8
`define GTME5_QUAD__CH1_RX_APT_CFG35_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG36    32'h000000d9
`define GTME5_QUAD__CH1_RX_APT_CFG36_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG37    32'h000000da
`define GTME5_QUAD__CH1_RX_APT_CFG37_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG38    32'h000000db
`define GTME5_QUAD__CH1_RX_APT_CFG38_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG39    32'h000000dc
`define GTME5_QUAD__CH1_RX_APT_CFG39_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG4    32'h000000dd
`define GTME5_QUAD__CH1_RX_APT_CFG4_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG40    32'h000000de
`define GTME5_QUAD__CH1_RX_APT_CFG40_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG41    32'h000000df
`define GTME5_QUAD__CH1_RX_APT_CFG41_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG42    32'h000000e0
`define GTME5_QUAD__CH1_RX_APT_CFG42_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG43    32'h000000e1
`define GTME5_QUAD__CH1_RX_APT_CFG43_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG44    32'h000000e2
`define GTME5_QUAD__CH1_RX_APT_CFG44_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG45    32'h000000e3
`define GTME5_QUAD__CH1_RX_APT_CFG45_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG46    32'h000000e4
`define GTME5_QUAD__CH1_RX_APT_CFG46_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG47    32'h000000e5
`define GTME5_QUAD__CH1_RX_APT_CFG47_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG48    32'h000000e6
`define GTME5_QUAD__CH1_RX_APT_CFG48_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG49    32'h000000e7
`define GTME5_QUAD__CH1_RX_APT_CFG49_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG5    32'h000000e8
`define GTME5_QUAD__CH1_RX_APT_CFG5_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG50    32'h000000e9
`define GTME5_QUAD__CH1_RX_APT_CFG50_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG51    32'h000000ea
`define GTME5_QUAD__CH1_RX_APT_CFG51_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG52    32'h000000eb
`define GTME5_QUAD__CH1_RX_APT_CFG52_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG53    32'h000000ec
`define GTME5_QUAD__CH1_RX_APT_CFG53_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG54    32'h000000ed
`define GTME5_QUAD__CH1_RX_APT_CFG54_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG55    32'h000000ee
`define GTME5_QUAD__CH1_RX_APT_CFG55_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG56    32'h000000ef
`define GTME5_QUAD__CH1_RX_APT_CFG56_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG57    32'h000000f0
`define GTME5_QUAD__CH1_RX_APT_CFG57_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG58    32'h000000f1
`define GTME5_QUAD__CH1_RX_APT_CFG58_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG6    32'h000000f2
`define GTME5_QUAD__CH1_RX_APT_CFG6_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG7    32'h000000f3
`define GTME5_QUAD__CH1_RX_APT_CFG7_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG8    32'h000000f4
`define GTME5_QUAD__CH1_RX_APT_CFG8_SZ 32

`define GTME5_QUAD__CH1_RX_APT_CFG9    32'h000000f5
`define GTME5_QUAD__CH1_RX_APT_CFG9_SZ 32

`define GTME5_QUAD__CH1_RX_CAL_CFG0    32'h000000f6
`define GTME5_QUAD__CH1_RX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_CAL_CFG1    32'h000000f7
`define GTME5_QUAD__CH1_RX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_CAL_CFG2    32'h000000f8
`define GTME5_QUAD__CH1_RX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG0    32'h000000f9
`define GTME5_QUAD__CH1_RX_CDR_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG1    32'h000000fa
`define GTME5_QUAD__CH1_RX_CDR_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG2    32'h000000fb
`define GTME5_QUAD__CH1_RX_CDR_CFG2_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG3    32'h000000fc
`define GTME5_QUAD__CH1_RX_CDR_CFG3_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG4    32'h000000fd
`define GTME5_QUAD__CH1_RX_CDR_CFG4_SZ 32

`define GTME5_QUAD__CH1_RX_CDR_CFG5    32'h000000fe
`define GTME5_QUAD__CH1_RX_CDR_CFG5_SZ 32

`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG0    32'h000000ff
`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG1    32'h00000100
`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG2    32'h00000101
`define GTME5_QUAD__CH1_RX_CTLE_ADC_CFG2_SZ 32

`define GTME5_QUAD__CH1_RX_CTLE_HF_CFG0    32'h00000102
`define GTME5_QUAD__CH1_RX_CTLE_HF_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_CTLE_HF_CFG1    32'h00000103
`define GTME5_QUAD__CH1_RX_CTLE_HF_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_DSP_CFG0    32'h00000104
`define GTME5_QUAD__CH1_RX_DSP_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_DSP_CFG1    32'h00000105
`define GTME5_QUAD__CH1_RX_DSP_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_MISC_CFG1    32'h00000106
`define GTME5_QUAD__CH1_RX_MISC_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_PAD_CFG0    32'h00000107
`define GTME5_QUAD__CH1_RX_PAD_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_PAD_CFG1    32'h00000108
`define GTME5_QUAD__CH1_RX_PAD_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_PCS_CFG0    32'h00000109
`define GTME5_QUAD__CH1_RX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_PCS_CFG1    32'h0000010a
`define GTME5_QUAD__CH1_RX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_RSV_CFG0    32'h0000010b
`define GTME5_QUAD__CH1_RX_RSV_CFG0_SZ 32

`define GTME5_QUAD__CH1_RX_RSV_CFG1    32'h0000010c
`define GTME5_QUAD__CH1_RX_RSV_CFG1_SZ 32

`define GTME5_QUAD__CH1_RX_SPARE_CFG0    32'h0000010d
`define GTME5_QUAD__CH1_RX_SPARE_CFG0_SZ 32

`define GTME5_QUAD__CH1_SIM_MODE    32'h0000010e
`define GTME5_QUAD__CH1_SIM_MODE_SZ 48

`define GTME5_QUAD__CH1_SIM_RECEIVER_DETECT_PASS    32'h0000010f
`define GTME5_QUAD__CH1_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTME5_QUAD__CH1_SIM_RESET_SPEEDUP    32'h00000110
`define GTME5_QUAD__CH1_SIM_RESET_SPEEDUP_SZ 40

`define GTME5_QUAD__CH1_TXOUTCLK_FREQ    32'h00000111
`define GTME5_QUAD__CH1_TXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH1_TXOUTCLK_REF_FREQ    32'h00000112
`define GTME5_QUAD__CH1_TXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH1_TXOUTCLK_REF_SOURCE    32'h00000113
`define GTME5_QUAD__CH1_TXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH1_TX_CAL_CFG0    32'h00000114
`define GTME5_QUAD__CH1_TX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH1_TX_CAL_CFG1    32'h00000115
`define GTME5_QUAD__CH1_TX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH1_TX_CAL_CFG2    32'h00000116
`define GTME5_QUAD__CH1_TX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH1_TX_CTRL_CFG0    32'h00000117
`define GTME5_QUAD__CH1_TX_CTRL_CFG0_SZ 32

`define GTME5_QUAD__CH1_TX_CTRL_CFG1    32'h00000118
`define GTME5_QUAD__CH1_TX_CTRL_CFG1_SZ 32

`define GTME5_QUAD__CH1_TX_CTRL_CFG2    32'h00000119
`define GTME5_QUAD__CH1_TX_CTRL_CFG2_SZ 32

`define GTME5_QUAD__CH1_TX_CTRL_CFG3    32'h0000011a
`define GTME5_QUAD__CH1_TX_CTRL_CFG3_SZ 32

`define GTME5_QUAD__CH1_TX_MISC_CFG0    32'h0000011b
`define GTME5_QUAD__CH1_TX_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG0    32'h0000011c
`define GTME5_QUAD__CH1_TX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG1    32'h0000011d
`define GTME5_QUAD__CH1_TX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG2    32'h0000011e
`define GTME5_QUAD__CH1_TX_PCS_CFG2_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG3    32'h0000011f
`define GTME5_QUAD__CH1_TX_PCS_CFG3_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG4    32'h00000120
`define GTME5_QUAD__CH1_TX_PCS_CFG4_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG5    32'h00000121
`define GTME5_QUAD__CH1_TX_PCS_CFG5_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG6    32'h00000122
`define GTME5_QUAD__CH1_TX_PCS_CFG6_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG7    32'h00000123
`define GTME5_QUAD__CH1_TX_PCS_CFG7_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG8    32'h00000124
`define GTME5_QUAD__CH1_TX_PCS_CFG8_SZ 32

`define GTME5_QUAD__CH1_TX_PCS_CFG9    32'h00000125
`define GTME5_QUAD__CH1_TX_PCS_CFG9_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG0    32'h00000126
`define GTME5_QUAD__CH2_CHCLK_CFG0_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG1    32'h00000127
`define GTME5_QUAD__CH2_CHCLK_CFG1_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG2    32'h00000128
`define GTME5_QUAD__CH2_CHCLK_CFG2_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG3    32'h00000129
`define GTME5_QUAD__CH2_CHCLK_CFG3_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG4    32'h0000012a
`define GTME5_QUAD__CH2_CHCLK_CFG4_SZ 32

`define GTME5_QUAD__CH2_CHCLK_CFG5    32'h0000012b
`define GTME5_QUAD__CH2_CHCLK_CFG5_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG0    32'h0000012c
`define GTME5_QUAD__CH2_EYESCAN_CFG0_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG1    32'h0000012d
`define GTME5_QUAD__CH2_EYESCAN_CFG1_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG2    32'h0000012e
`define GTME5_QUAD__CH2_EYESCAN_CFG2_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG3    32'h0000012f
`define GTME5_QUAD__CH2_EYESCAN_CFG3_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG4    32'h00000130
`define GTME5_QUAD__CH2_EYESCAN_CFG4_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG5    32'h00000131
`define GTME5_QUAD__CH2_EYESCAN_CFG5_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG6    32'h00000132
`define GTME5_QUAD__CH2_EYESCAN_CFG6_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG7    32'h00000133
`define GTME5_QUAD__CH2_EYESCAN_CFG7_SZ 32

`define GTME5_QUAD__CH2_EYESCAN_CFG8    32'h00000134
`define GTME5_QUAD__CH2_EYESCAN_CFG8_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG0    32'h00000135
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG0_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG1    32'h00000136
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG1_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG2    32'h00000137
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG2_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG3    32'h00000138
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG3_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG4    32'h00000139
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG4_SZ 32

`define GTME5_QUAD__CH2_FABRIC_INTF_CFG5    32'h0000013a
`define GTME5_QUAD__CH2_FABRIC_INTF_CFG5_SZ 32

`define GTME5_QUAD__CH2_INSTANTIATED    32'h0000013b
`define GTME5_QUAD__CH2_INSTANTIATED_SZ 1

`define GTME5_QUAD__CH2_MONITOR_CFG0    32'h0000013c
`define GTME5_QUAD__CH2_MONITOR_CFG0_SZ 32

`define GTME5_QUAD__CH2_PMA_MISC_CFG0    32'h0000013d
`define GTME5_QUAD__CH2_PMA_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH2_RESET_BYP_HDSHK_CFG    32'h0000013e
`define GTME5_QUAD__CH2_RESET_BYP_HDSHK_CFG_SZ 32

`define GTME5_QUAD__CH2_RESET_CFG    32'h0000013f
`define GTME5_QUAD__CH2_RESET_CFG_SZ 32

`define GTME5_QUAD__CH2_RESET_LOOPER_ID_CFG    32'h00000140
`define GTME5_QUAD__CH2_RESET_LOOPER_ID_CFG_SZ 32

`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG0    32'h00000141
`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG0_SZ 32

`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG1    32'h00000142
`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG1_SZ 32

`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG2    32'h00000143
`define GTME5_QUAD__CH2_RESET_LOOP_ID_CFG2_SZ 32

`define GTME5_QUAD__CH2_RESET_TIME_CFG0    32'h00000144
`define GTME5_QUAD__CH2_RESET_TIME_CFG0_SZ 32

`define GTME5_QUAD__CH2_RESET_TIME_CFG1    32'h00000145
`define GTME5_QUAD__CH2_RESET_TIME_CFG1_SZ 32

`define GTME5_QUAD__CH2_RESET_TIME_CFG2    32'h00000146
`define GTME5_QUAD__CH2_RESET_TIME_CFG2_SZ 32

`define GTME5_QUAD__CH2_RESET_TIME_CFG3    32'h00000147
`define GTME5_QUAD__CH2_RESET_TIME_CFG3_SZ 32

`define GTME5_QUAD__CH2_RXOUTCLK_FREQ    32'h00000148
`define GTME5_QUAD__CH2_RXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH2_RXOUTCLK_REF_FREQ    32'h00000149
`define GTME5_QUAD__CH2_RXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH2_RXOUTCLK_REF_SOURCE    32'h0000014a
`define GTME5_QUAD__CH2_RXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH2_RX_APT_CFG0    32'h0000014b
`define GTME5_QUAD__CH2_RX_APT_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG1    32'h0000014c
`define GTME5_QUAD__CH2_RX_APT_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG10    32'h0000014d
`define GTME5_QUAD__CH2_RX_APT_CFG10_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG11    32'h0000014e
`define GTME5_QUAD__CH2_RX_APT_CFG11_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG12    32'h0000014f
`define GTME5_QUAD__CH2_RX_APT_CFG12_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG13    32'h00000150
`define GTME5_QUAD__CH2_RX_APT_CFG13_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG14    32'h00000151
`define GTME5_QUAD__CH2_RX_APT_CFG14_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG15    32'h00000152
`define GTME5_QUAD__CH2_RX_APT_CFG15_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG16    32'h00000153
`define GTME5_QUAD__CH2_RX_APT_CFG16_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG17    32'h00000154
`define GTME5_QUAD__CH2_RX_APT_CFG17_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG18    32'h00000155
`define GTME5_QUAD__CH2_RX_APT_CFG18_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG19    32'h00000156
`define GTME5_QUAD__CH2_RX_APT_CFG19_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG2    32'h00000157
`define GTME5_QUAD__CH2_RX_APT_CFG2_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG20    32'h00000158
`define GTME5_QUAD__CH2_RX_APT_CFG20_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG21    32'h00000159
`define GTME5_QUAD__CH2_RX_APT_CFG21_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG22    32'h0000015a
`define GTME5_QUAD__CH2_RX_APT_CFG22_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG23    32'h0000015b
`define GTME5_QUAD__CH2_RX_APT_CFG23_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG24    32'h0000015c
`define GTME5_QUAD__CH2_RX_APT_CFG24_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG25    32'h0000015d
`define GTME5_QUAD__CH2_RX_APT_CFG25_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG26    32'h0000015e
`define GTME5_QUAD__CH2_RX_APT_CFG26_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG27    32'h0000015f
`define GTME5_QUAD__CH2_RX_APT_CFG27_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG28    32'h00000160
`define GTME5_QUAD__CH2_RX_APT_CFG28_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG29    32'h00000161
`define GTME5_QUAD__CH2_RX_APT_CFG29_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG3    32'h00000162
`define GTME5_QUAD__CH2_RX_APT_CFG3_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG30    32'h00000163
`define GTME5_QUAD__CH2_RX_APT_CFG30_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG31    32'h00000164
`define GTME5_QUAD__CH2_RX_APT_CFG31_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG32    32'h00000165
`define GTME5_QUAD__CH2_RX_APT_CFG32_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG33    32'h00000166
`define GTME5_QUAD__CH2_RX_APT_CFG33_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG34    32'h00000167
`define GTME5_QUAD__CH2_RX_APT_CFG34_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG35    32'h00000168
`define GTME5_QUAD__CH2_RX_APT_CFG35_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG36    32'h00000169
`define GTME5_QUAD__CH2_RX_APT_CFG36_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG37    32'h0000016a
`define GTME5_QUAD__CH2_RX_APT_CFG37_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG38    32'h0000016b
`define GTME5_QUAD__CH2_RX_APT_CFG38_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG39    32'h0000016c
`define GTME5_QUAD__CH2_RX_APT_CFG39_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG4    32'h0000016d
`define GTME5_QUAD__CH2_RX_APT_CFG4_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG40    32'h0000016e
`define GTME5_QUAD__CH2_RX_APT_CFG40_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG41    32'h0000016f
`define GTME5_QUAD__CH2_RX_APT_CFG41_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG42    32'h00000170
`define GTME5_QUAD__CH2_RX_APT_CFG42_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG43    32'h00000171
`define GTME5_QUAD__CH2_RX_APT_CFG43_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG44    32'h00000172
`define GTME5_QUAD__CH2_RX_APT_CFG44_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG45    32'h00000173
`define GTME5_QUAD__CH2_RX_APT_CFG45_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG46    32'h00000174
`define GTME5_QUAD__CH2_RX_APT_CFG46_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG47    32'h00000175
`define GTME5_QUAD__CH2_RX_APT_CFG47_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG48    32'h00000176
`define GTME5_QUAD__CH2_RX_APT_CFG48_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG49    32'h00000177
`define GTME5_QUAD__CH2_RX_APT_CFG49_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG5    32'h00000178
`define GTME5_QUAD__CH2_RX_APT_CFG5_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG50    32'h00000179
`define GTME5_QUAD__CH2_RX_APT_CFG50_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG51    32'h0000017a
`define GTME5_QUAD__CH2_RX_APT_CFG51_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG52    32'h0000017b
`define GTME5_QUAD__CH2_RX_APT_CFG52_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG53    32'h0000017c
`define GTME5_QUAD__CH2_RX_APT_CFG53_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG54    32'h0000017d
`define GTME5_QUAD__CH2_RX_APT_CFG54_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG55    32'h0000017e
`define GTME5_QUAD__CH2_RX_APT_CFG55_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG56    32'h0000017f
`define GTME5_QUAD__CH2_RX_APT_CFG56_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG57    32'h00000180
`define GTME5_QUAD__CH2_RX_APT_CFG57_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG58    32'h00000181
`define GTME5_QUAD__CH2_RX_APT_CFG58_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG6    32'h00000182
`define GTME5_QUAD__CH2_RX_APT_CFG6_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG7    32'h00000183
`define GTME5_QUAD__CH2_RX_APT_CFG7_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG8    32'h00000184
`define GTME5_QUAD__CH2_RX_APT_CFG8_SZ 32

`define GTME5_QUAD__CH2_RX_APT_CFG9    32'h00000185
`define GTME5_QUAD__CH2_RX_APT_CFG9_SZ 32

`define GTME5_QUAD__CH2_RX_CAL_CFG0    32'h00000186
`define GTME5_QUAD__CH2_RX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_CAL_CFG1    32'h00000187
`define GTME5_QUAD__CH2_RX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_CAL_CFG2    32'h00000188
`define GTME5_QUAD__CH2_RX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG0    32'h00000189
`define GTME5_QUAD__CH2_RX_CDR_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG1    32'h0000018a
`define GTME5_QUAD__CH2_RX_CDR_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG2    32'h0000018b
`define GTME5_QUAD__CH2_RX_CDR_CFG2_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG3    32'h0000018c
`define GTME5_QUAD__CH2_RX_CDR_CFG3_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG4    32'h0000018d
`define GTME5_QUAD__CH2_RX_CDR_CFG4_SZ 32

`define GTME5_QUAD__CH2_RX_CDR_CFG5    32'h0000018e
`define GTME5_QUAD__CH2_RX_CDR_CFG5_SZ 32

`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG0    32'h0000018f
`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG1    32'h00000190
`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG2    32'h00000191
`define GTME5_QUAD__CH2_RX_CTLE_ADC_CFG2_SZ 32

`define GTME5_QUAD__CH2_RX_CTLE_HF_CFG0    32'h00000192
`define GTME5_QUAD__CH2_RX_CTLE_HF_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_CTLE_HF_CFG1    32'h00000193
`define GTME5_QUAD__CH2_RX_CTLE_HF_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_DSP_CFG0    32'h00000194
`define GTME5_QUAD__CH2_RX_DSP_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_DSP_CFG1    32'h00000195
`define GTME5_QUAD__CH2_RX_DSP_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_MISC_CFG1    32'h00000196
`define GTME5_QUAD__CH2_RX_MISC_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_PAD_CFG0    32'h00000197
`define GTME5_QUAD__CH2_RX_PAD_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_PAD_CFG1    32'h00000198
`define GTME5_QUAD__CH2_RX_PAD_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_PCS_CFG0    32'h00000199
`define GTME5_QUAD__CH2_RX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_PCS_CFG1    32'h0000019a
`define GTME5_QUAD__CH2_RX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_RSV_CFG0    32'h0000019b
`define GTME5_QUAD__CH2_RX_RSV_CFG0_SZ 32

`define GTME5_QUAD__CH2_RX_RSV_CFG1    32'h0000019c
`define GTME5_QUAD__CH2_RX_RSV_CFG1_SZ 32

`define GTME5_QUAD__CH2_RX_SPARE_CFG0    32'h0000019d
`define GTME5_QUAD__CH2_RX_SPARE_CFG0_SZ 32

`define GTME5_QUAD__CH2_SIM_MODE    32'h0000019e
`define GTME5_QUAD__CH2_SIM_MODE_SZ 48

`define GTME5_QUAD__CH2_SIM_RECEIVER_DETECT_PASS    32'h0000019f
`define GTME5_QUAD__CH2_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTME5_QUAD__CH2_SIM_RESET_SPEEDUP    32'h000001a0
`define GTME5_QUAD__CH2_SIM_RESET_SPEEDUP_SZ 40

`define GTME5_QUAD__CH2_TXOUTCLK_FREQ    32'h000001a1
`define GTME5_QUAD__CH2_TXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH2_TXOUTCLK_REF_FREQ    32'h000001a2
`define GTME5_QUAD__CH2_TXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH2_TXOUTCLK_REF_SOURCE    32'h000001a3
`define GTME5_QUAD__CH2_TXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH2_TX_CAL_CFG0    32'h000001a4
`define GTME5_QUAD__CH2_TX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH2_TX_CAL_CFG1    32'h000001a5
`define GTME5_QUAD__CH2_TX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH2_TX_CAL_CFG2    32'h000001a6
`define GTME5_QUAD__CH2_TX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH2_TX_CTRL_CFG0    32'h000001a7
`define GTME5_QUAD__CH2_TX_CTRL_CFG0_SZ 32

`define GTME5_QUAD__CH2_TX_CTRL_CFG1    32'h000001a8
`define GTME5_QUAD__CH2_TX_CTRL_CFG1_SZ 32

`define GTME5_QUAD__CH2_TX_CTRL_CFG2    32'h000001a9
`define GTME5_QUAD__CH2_TX_CTRL_CFG2_SZ 32

`define GTME5_QUAD__CH2_TX_CTRL_CFG3    32'h000001aa
`define GTME5_QUAD__CH2_TX_CTRL_CFG3_SZ 32

`define GTME5_QUAD__CH2_TX_MISC_CFG0    32'h000001ab
`define GTME5_QUAD__CH2_TX_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG0    32'h000001ac
`define GTME5_QUAD__CH2_TX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG1    32'h000001ad
`define GTME5_QUAD__CH2_TX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG2    32'h000001ae
`define GTME5_QUAD__CH2_TX_PCS_CFG2_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG3    32'h000001af
`define GTME5_QUAD__CH2_TX_PCS_CFG3_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG4    32'h000001b0
`define GTME5_QUAD__CH2_TX_PCS_CFG4_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG5    32'h000001b1
`define GTME5_QUAD__CH2_TX_PCS_CFG5_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG6    32'h000001b2
`define GTME5_QUAD__CH2_TX_PCS_CFG6_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG7    32'h000001b3
`define GTME5_QUAD__CH2_TX_PCS_CFG7_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG8    32'h000001b4
`define GTME5_QUAD__CH2_TX_PCS_CFG8_SZ 32

`define GTME5_QUAD__CH2_TX_PCS_CFG9    32'h000001b5
`define GTME5_QUAD__CH2_TX_PCS_CFG9_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG0    32'h000001b6
`define GTME5_QUAD__CH3_CHCLK_CFG0_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG1    32'h000001b7
`define GTME5_QUAD__CH3_CHCLK_CFG1_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG2    32'h000001b8
`define GTME5_QUAD__CH3_CHCLK_CFG2_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG3    32'h000001b9
`define GTME5_QUAD__CH3_CHCLK_CFG3_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG4    32'h000001ba
`define GTME5_QUAD__CH3_CHCLK_CFG4_SZ 32

`define GTME5_QUAD__CH3_CHCLK_CFG5    32'h000001bb
`define GTME5_QUAD__CH3_CHCLK_CFG5_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG0    32'h000001bc
`define GTME5_QUAD__CH3_EYESCAN_CFG0_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG1    32'h000001bd
`define GTME5_QUAD__CH3_EYESCAN_CFG1_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG2    32'h000001be
`define GTME5_QUAD__CH3_EYESCAN_CFG2_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG3    32'h000001bf
`define GTME5_QUAD__CH3_EYESCAN_CFG3_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG4    32'h000001c0
`define GTME5_QUAD__CH3_EYESCAN_CFG4_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG5    32'h000001c1
`define GTME5_QUAD__CH3_EYESCAN_CFG5_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG6    32'h000001c2
`define GTME5_QUAD__CH3_EYESCAN_CFG6_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG7    32'h000001c3
`define GTME5_QUAD__CH3_EYESCAN_CFG7_SZ 32

`define GTME5_QUAD__CH3_EYESCAN_CFG8    32'h000001c4
`define GTME5_QUAD__CH3_EYESCAN_CFG8_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG0    32'h000001c5
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG0_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG1    32'h000001c6
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG1_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG2    32'h000001c7
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG2_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG3    32'h000001c8
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG3_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG4    32'h000001c9
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG4_SZ 32

`define GTME5_QUAD__CH3_FABRIC_INTF_CFG5    32'h000001ca
`define GTME5_QUAD__CH3_FABRIC_INTF_CFG5_SZ 32

`define GTME5_QUAD__CH3_INSTANTIATED    32'h000001cb
`define GTME5_QUAD__CH3_INSTANTIATED_SZ 1

`define GTME5_QUAD__CH3_MONITOR_CFG0    32'h000001cc
`define GTME5_QUAD__CH3_MONITOR_CFG0_SZ 32

`define GTME5_QUAD__CH3_PMA_MISC_CFG0    32'h000001cd
`define GTME5_QUAD__CH3_PMA_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH3_RESET_BYP_HDSHK_CFG    32'h000001ce
`define GTME5_QUAD__CH3_RESET_BYP_HDSHK_CFG_SZ 32

`define GTME5_QUAD__CH3_RESET_CFG    32'h000001cf
`define GTME5_QUAD__CH3_RESET_CFG_SZ 32

`define GTME5_QUAD__CH3_RESET_LOOPER_ID_CFG    32'h000001d0
`define GTME5_QUAD__CH3_RESET_LOOPER_ID_CFG_SZ 32

`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG0    32'h000001d1
`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG0_SZ 32

`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG1    32'h000001d2
`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG1_SZ 32

`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG2    32'h000001d3
`define GTME5_QUAD__CH3_RESET_LOOP_ID_CFG2_SZ 32

`define GTME5_QUAD__CH3_RESET_TIME_CFG0    32'h000001d4
`define GTME5_QUAD__CH3_RESET_TIME_CFG0_SZ 32

`define GTME5_QUAD__CH3_RESET_TIME_CFG1    32'h000001d5
`define GTME5_QUAD__CH3_RESET_TIME_CFG1_SZ 32

`define GTME5_QUAD__CH3_RESET_TIME_CFG2    32'h000001d6
`define GTME5_QUAD__CH3_RESET_TIME_CFG2_SZ 32

`define GTME5_QUAD__CH3_RESET_TIME_CFG3    32'h000001d7
`define GTME5_QUAD__CH3_RESET_TIME_CFG3_SZ 32

`define GTME5_QUAD__CH3_RXOUTCLK_FREQ    32'h000001d8
`define GTME5_QUAD__CH3_RXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH3_RXOUTCLK_REF_FREQ    32'h000001d9
`define GTME5_QUAD__CH3_RXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH3_RXOUTCLK_REF_SOURCE    32'h000001da
`define GTME5_QUAD__CH3_RXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH3_RX_APT_CFG0    32'h000001db
`define GTME5_QUAD__CH3_RX_APT_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG1    32'h000001dc
`define GTME5_QUAD__CH3_RX_APT_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG10    32'h000001dd
`define GTME5_QUAD__CH3_RX_APT_CFG10_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG11    32'h000001de
`define GTME5_QUAD__CH3_RX_APT_CFG11_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG12    32'h000001df
`define GTME5_QUAD__CH3_RX_APT_CFG12_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG13    32'h000001e0
`define GTME5_QUAD__CH3_RX_APT_CFG13_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG14    32'h000001e1
`define GTME5_QUAD__CH3_RX_APT_CFG14_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG15    32'h000001e2
`define GTME5_QUAD__CH3_RX_APT_CFG15_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG16    32'h000001e3
`define GTME5_QUAD__CH3_RX_APT_CFG16_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG17    32'h000001e4
`define GTME5_QUAD__CH3_RX_APT_CFG17_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG18    32'h000001e5
`define GTME5_QUAD__CH3_RX_APT_CFG18_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG19    32'h000001e6
`define GTME5_QUAD__CH3_RX_APT_CFG19_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG2    32'h000001e7
`define GTME5_QUAD__CH3_RX_APT_CFG2_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG20    32'h000001e8
`define GTME5_QUAD__CH3_RX_APT_CFG20_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG21    32'h000001e9
`define GTME5_QUAD__CH3_RX_APT_CFG21_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG22    32'h000001ea
`define GTME5_QUAD__CH3_RX_APT_CFG22_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG23    32'h000001eb
`define GTME5_QUAD__CH3_RX_APT_CFG23_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG24    32'h000001ec
`define GTME5_QUAD__CH3_RX_APT_CFG24_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG25    32'h000001ed
`define GTME5_QUAD__CH3_RX_APT_CFG25_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG26    32'h000001ee
`define GTME5_QUAD__CH3_RX_APT_CFG26_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG27    32'h000001ef
`define GTME5_QUAD__CH3_RX_APT_CFG27_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG28    32'h000001f0
`define GTME5_QUAD__CH3_RX_APT_CFG28_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG29    32'h000001f1
`define GTME5_QUAD__CH3_RX_APT_CFG29_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG3    32'h000001f2
`define GTME5_QUAD__CH3_RX_APT_CFG3_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG30    32'h000001f3
`define GTME5_QUAD__CH3_RX_APT_CFG30_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG31    32'h000001f4
`define GTME5_QUAD__CH3_RX_APT_CFG31_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG32    32'h000001f5
`define GTME5_QUAD__CH3_RX_APT_CFG32_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG33    32'h000001f6
`define GTME5_QUAD__CH3_RX_APT_CFG33_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG34    32'h000001f7
`define GTME5_QUAD__CH3_RX_APT_CFG34_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG35    32'h000001f8
`define GTME5_QUAD__CH3_RX_APT_CFG35_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG36    32'h000001f9
`define GTME5_QUAD__CH3_RX_APT_CFG36_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG37    32'h000001fa
`define GTME5_QUAD__CH3_RX_APT_CFG37_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG38    32'h000001fb
`define GTME5_QUAD__CH3_RX_APT_CFG38_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG39    32'h000001fc
`define GTME5_QUAD__CH3_RX_APT_CFG39_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG4    32'h000001fd
`define GTME5_QUAD__CH3_RX_APT_CFG4_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG40    32'h000001fe
`define GTME5_QUAD__CH3_RX_APT_CFG40_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG41    32'h000001ff
`define GTME5_QUAD__CH3_RX_APT_CFG41_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG42    32'h00000200
`define GTME5_QUAD__CH3_RX_APT_CFG42_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG43    32'h00000201
`define GTME5_QUAD__CH3_RX_APT_CFG43_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG44    32'h00000202
`define GTME5_QUAD__CH3_RX_APT_CFG44_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG45    32'h00000203
`define GTME5_QUAD__CH3_RX_APT_CFG45_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG46    32'h00000204
`define GTME5_QUAD__CH3_RX_APT_CFG46_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG47    32'h00000205
`define GTME5_QUAD__CH3_RX_APT_CFG47_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG48    32'h00000206
`define GTME5_QUAD__CH3_RX_APT_CFG48_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG49    32'h00000207
`define GTME5_QUAD__CH3_RX_APT_CFG49_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG5    32'h00000208
`define GTME5_QUAD__CH3_RX_APT_CFG5_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG50    32'h00000209
`define GTME5_QUAD__CH3_RX_APT_CFG50_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG51    32'h0000020a
`define GTME5_QUAD__CH3_RX_APT_CFG51_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG52    32'h0000020b
`define GTME5_QUAD__CH3_RX_APT_CFG52_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG53    32'h0000020c
`define GTME5_QUAD__CH3_RX_APT_CFG53_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG54    32'h0000020d
`define GTME5_QUAD__CH3_RX_APT_CFG54_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG55    32'h0000020e
`define GTME5_QUAD__CH3_RX_APT_CFG55_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG56    32'h0000020f
`define GTME5_QUAD__CH3_RX_APT_CFG56_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG57    32'h00000210
`define GTME5_QUAD__CH3_RX_APT_CFG57_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG58    32'h00000211
`define GTME5_QUAD__CH3_RX_APT_CFG58_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG6    32'h00000212
`define GTME5_QUAD__CH3_RX_APT_CFG6_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG7    32'h00000213
`define GTME5_QUAD__CH3_RX_APT_CFG7_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG8    32'h00000214
`define GTME5_QUAD__CH3_RX_APT_CFG8_SZ 32

`define GTME5_QUAD__CH3_RX_APT_CFG9    32'h00000215
`define GTME5_QUAD__CH3_RX_APT_CFG9_SZ 32

`define GTME5_QUAD__CH3_RX_CAL_CFG0    32'h00000216
`define GTME5_QUAD__CH3_RX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_CAL_CFG1    32'h00000217
`define GTME5_QUAD__CH3_RX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_CAL_CFG2    32'h00000218
`define GTME5_QUAD__CH3_RX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG0    32'h00000219
`define GTME5_QUAD__CH3_RX_CDR_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG1    32'h0000021a
`define GTME5_QUAD__CH3_RX_CDR_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG2    32'h0000021b
`define GTME5_QUAD__CH3_RX_CDR_CFG2_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG3    32'h0000021c
`define GTME5_QUAD__CH3_RX_CDR_CFG3_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG4    32'h0000021d
`define GTME5_QUAD__CH3_RX_CDR_CFG4_SZ 32

`define GTME5_QUAD__CH3_RX_CDR_CFG5    32'h0000021e
`define GTME5_QUAD__CH3_RX_CDR_CFG5_SZ 32

`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG0    32'h0000021f
`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG1    32'h00000220
`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG2    32'h00000221
`define GTME5_QUAD__CH3_RX_CTLE_ADC_CFG2_SZ 32

`define GTME5_QUAD__CH3_RX_CTLE_HF_CFG0    32'h00000222
`define GTME5_QUAD__CH3_RX_CTLE_HF_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_CTLE_HF_CFG1    32'h00000223
`define GTME5_QUAD__CH3_RX_CTLE_HF_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_DSP_CFG0    32'h00000224
`define GTME5_QUAD__CH3_RX_DSP_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_DSP_CFG1    32'h00000225
`define GTME5_QUAD__CH3_RX_DSP_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_MISC_CFG1    32'h00000226
`define GTME5_QUAD__CH3_RX_MISC_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_PAD_CFG0    32'h00000227
`define GTME5_QUAD__CH3_RX_PAD_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_PAD_CFG1    32'h00000228
`define GTME5_QUAD__CH3_RX_PAD_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_PCS_CFG0    32'h00000229
`define GTME5_QUAD__CH3_RX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_PCS_CFG1    32'h0000022a
`define GTME5_QUAD__CH3_RX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_RSV_CFG0    32'h0000022b
`define GTME5_QUAD__CH3_RX_RSV_CFG0_SZ 32

`define GTME5_QUAD__CH3_RX_RSV_CFG1    32'h0000022c
`define GTME5_QUAD__CH3_RX_RSV_CFG1_SZ 32

`define GTME5_QUAD__CH3_RX_SPARE_CFG0    32'h0000022d
`define GTME5_QUAD__CH3_RX_SPARE_CFG0_SZ 32

`define GTME5_QUAD__CH3_SIM_MODE    32'h0000022e
`define GTME5_QUAD__CH3_SIM_MODE_SZ 48

`define GTME5_QUAD__CH3_SIM_RECEIVER_DETECT_PASS    32'h0000022f
`define GTME5_QUAD__CH3_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTME5_QUAD__CH3_SIM_RESET_SPEEDUP    32'h00000230
`define GTME5_QUAD__CH3_SIM_RESET_SPEEDUP_SZ 40

`define GTME5_QUAD__CH3_TXOUTCLK_FREQ    32'h00000231
`define GTME5_QUAD__CH3_TXOUTCLK_FREQ_SZ 64

`define GTME5_QUAD__CH3_TXOUTCLK_REF_FREQ    32'h00000232
`define GTME5_QUAD__CH3_TXOUTCLK_REF_FREQ_SZ 64

`define GTME5_QUAD__CH3_TXOUTCLK_REF_SOURCE    32'h00000233
`define GTME5_QUAD__CH3_TXOUTCLK_REF_SOURCE_SZ 192

`define GTME5_QUAD__CH3_TX_CAL_CFG0    32'h00000234
`define GTME5_QUAD__CH3_TX_CAL_CFG0_SZ 32

`define GTME5_QUAD__CH3_TX_CAL_CFG1    32'h00000235
`define GTME5_QUAD__CH3_TX_CAL_CFG1_SZ 32

`define GTME5_QUAD__CH3_TX_CAL_CFG2    32'h00000236
`define GTME5_QUAD__CH3_TX_CAL_CFG2_SZ 32

`define GTME5_QUAD__CH3_TX_CTRL_CFG0    32'h00000237
`define GTME5_QUAD__CH3_TX_CTRL_CFG0_SZ 32

`define GTME5_QUAD__CH3_TX_CTRL_CFG1    32'h00000238
`define GTME5_QUAD__CH3_TX_CTRL_CFG1_SZ 32

`define GTME5_QUAD__CH3_TX_CTRL_CFG2    32'h00000239
`define GTME5_QUAD__CH3_TX_CTRL_CFG2_SZ 32

`define GTME5_QUAD__CH3_TX_CTRL_CFG3    32'h0000023a
`define GTME5_QUAD__CH3_TX_CTRL_CFG3_SZ 32

`define GTME5_QUAD__CH3_TX_MISC_CFG0    32'h0000023b
`define GTME5_QUAD__CH3_TX_MISC_CFG0_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG0    32'h0000023c
`define GTME5_QUAD__CH3_TX_PCS_CFG0_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG1    32'h0000023d
`define GTME5_QUAD__CH3_TX_PCS_CFG1_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG2    32'h0000023e
`define GTME5_QUAD__CH3_TX_PCS_CFG2_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG3    32'h0000023f
`define GTME5_QUAD__CH3_TX_PCS_CFG3_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG4    32'h00000240
`define GTME5_QUAD__CH3_TX_PCS_CFG4_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG5    32'h00000241
`define GTME5_QUAD__CH3_TX_PCS_CFG5_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG6    32'h00000242
`define GTME5_QUAD__CH3_TX_PCS_CFG6_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG7    32'h00000243
`define GTME5_QUAD__CH3_TX_PCS_CFG7_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG8    32'h00000244
`define GTME5_QUAD__CH3_TX_PCS_CFG8_SZ 32

`define GTME5_QUAD__CH3_TX_PCS_CFG9    32'h00000245
`define GTME5_QUAD__CH3_TX_PCS_CFG9_SZ 32

`define GTME5_QUAD__CHANNEL_CONNECTIVITY    32'h00000246
`define GTME5_QUAD__CHANNEL_CONNECTIVITY_SZ 32

`define GTME5_QUAD__CTRL_RSV_CFG0    32'h00000247
`define GTME5_QUAD__CTRL_RSV_CFG0_SZ 32

`define GTME5_QUAD__CTRL_RSV_CFG1    32'h00000248
`define GTME5_QUAD__CTRL_RSV_CFG1_SZ 32

`define GTME5_QUAD__HS0_LCPLL_IPS_PIN_EN    32'h00000249
`define GTME5_QUAD__HS0_LCPLL_IPS_PIN_EN_SZ 1

`define GTME5_QUAD__HS0_LCPLL_IPS_REFCLK_SEL    32'h0000024a
`define GTME5_QUAD__HS0_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP0    32'h0000024b
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP0_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP1    32'h0000024c
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP1_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP2    32'h0000024d
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP2_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP3    32'h0000024e
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP3_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP4    32'h0000024f
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP4_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP5    32'h00000250
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP5_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP6    32'h00000251
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP6_SZ 3

`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP7    32'h00000252
`define GTME5_QUAD__HS0_LCPLL_REFCLK_MAP7_SZ 3

`define GTME5_QUAD__HS1_LCPLL_IPS_PIN_EN    32'h00000253
`define GTME5_QUAD__HS1_LCPLL_IPS_PIN_EN_SZ 1

`define GTME5_QUAD__HS1_LCPLL_IPS_REFCLK_SEL    32'h00000254
`define GTME5_QUAD__HS1_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP0    32'h00000255
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP0_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP1    32'h00000256
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP1_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP2    32'h00000257
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP2_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP3    32'h00000258
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP3_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP4    32'h00000259
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP4_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP5    32'h0000025a
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP5_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP6    32'h0000025b
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP6_SZ 3

`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP7    32'h0000025c
`define GTME5_QUAD__HS1_LCPLL_REFCLK_MAP7_SZ 3

`define GTME5_QUAD__HSCLK0_HSDIST_CFG    32'h0000025d
`define GTME5_QUAD__HSCLK0_HSDIST_CFG_SZ 32

`define GTME5_QUAD__HSCLK0_INSTANTIATED    32'h0000025e
`define GTME5_QUAD__HSCLK0_INSTANTIATED_SZ 1

`define GTME5_QUAD__HSCLK0_LCPLL_CFG0    32'h0000025f
`define GTME5_QUAD__HSCLK0_LCPLL_CFG0_SZ 32

`define GTME5_QUAD__HSCLK0_LCPLL_CFG1    32'h00000260
`define GTME5_QUAD__HSCLK0_LCPLL_CFG1_SZ 32

`define GTME5_QUAD__HSCLK0_LCPLL_CFG2    32'h00000261
`define GTME5_QUAD__HSCLK0_LCPLL_CFG2_SZ 32

`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG0    32'h00000262
`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG0_SZ 32

`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG1    32'h00000263
`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG1_SZ 32

`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG2    32'h00000264
`define GTME5_QUAD__HSCLK0_LCPLL_LGC_CFG2_SZ 32

`define GTME5_QUAD__HSCLK0_RXRECCLK_SEL    32'h00000265
`define GTME5_QUAD__HSCLK0_RXRECCLK_SEL_SZ 2

`define GTME5_QUAD__HSCLK1_HSDIST_CFG    32'h00000266
`define GTME5_QUAD__HSCLK1_HSDIST_CFG_SZ 32

`define GTME5_QUAD__HSCLK1_INSTANTIATED    32'h00000267
`define GTME5_QUAD__HSCLK1_INSTANTIATED_SZ 1

`define GTME5_QUAD__HSCLK1_LCPLL_CFG0    32'h00000268
`define GTME5_QUAD__HSCLK1_LCPLL_CFG0_SZ 32

`define GTME5_QUAD__HSCLK1_LCPLL_CFG1    32'h00000269
`define GTME5_QUAD__HSCLK1_LCPLL_CFG1_SZ 32

`define GTME5_QUAD__HSCLK1_LCPLL_CFG2    32'h0000026a
`define GTME5_QUAD__HSCLK1_LCPLL_CFG2_SZ 32

`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG0    32'h0000026b
`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG0_SZ 32

`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG1    32'h0000026c
`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG1_SZ 32

`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG2    32'h0000026d
`define GTME5_QUAD__HSCLK1_LCPLL_LGC_CFG2_SZ 32

`define GTME5_QUAD__HSCLK1_RXRECCLK_SEL    32'h0000026e
`define GTME5_QUAD__HSCLK1_RXRECCLK_SEL_SZ 2

`define GTME5_QUAD__MEMORY_INIT_FILE    32'h0000026f
`define GTME5_QUAD__MEMORY_INIT_FILE_SZ 32

`define GTME5_QUAD__MST_RESET_CFG    32'h00000270
`define GTME5_QUAD__MST_RESET_CFG_SZ 32

`define GTME5_QUAD__PIN_CFG0    32'h00000271
`define GTME5_QUAD__PIN_CFG0_SZ 32

`define GTME5_QUAD__POR_CFG    32'h00000272
`define GTME5_QUAD__POR_CFG_SZ 32

`define GTME5_QUAD__QUAD_INSTANTIATED    32'h00000273
`define GTME5_QUAD__QUAD_INSTANTIATED_SZ 1

`define GTME5_QUAD__QUAD_SIM_MODE    32'h00000274
`define GTME5_QUAD__QUAD_SIM_MODE_SZ 48

`define GTME5_QUAD__QUAD_SIM_RESET_SPEEDUP    32'h00000275
`define GTME5_QUAD__QUAD_SIM_RESET_SPEEDUP_SZ 40

`define GTME5_QUAD__RCALBG0_CFG0    32'h00000276
`define GTME5_QUAD__RCALBG0_CFG0_SZ 32

`define GTME5_QUAD__RCALBG0_CFG1    32'h00000277
`define GTME5_QUAD__RCALBG0_CFG1_SZ 32

`define GTME5_QUAD__RCALBG0_CFG2    32'h00000278
`define GTME5_QUAD__RCALBG0_CFG2_SZ 32

`define GTME5_QUAD__RCALBG0_CFG3    32'h00000279
`define GTME5_QUAD__RCALBG0_CFG3_SZ 32

`define GTME5_QUAD__RCALBG0_CFG4    32'h0000027a
`define GTME5_QUAD__RCALBG0_CFG4_SZ 32

`define GTME5_QUAD__RCALBG0_CFG5    32'h0000027b
`define GTME5_QUAD__RCALBG0_CFG5_SZ 32

`define GTME5_QUAD__RCALBG1_CFG0    32'h0000027c
`define GTME5_QUAD__RCALBG1_CFG0_SZ 32

`define GTME5_QUAD__RCALBG1_CFG1    32'h0000027d
`define GTME5_QUAD__RCALBG1_CFG1_SZ 32

`define GTME5_QUAD__RCALBG1_CFG2    32'h0000027e
`define GTME5_QUAD__RCALBG1_CFG2_SZ 32

`define GTME5_QUAD__RCALBG1_CFG3    32'h0000027f
`define GTME5_QUAD__RCALBG1_CFG3_SZ 32

`define GTME5_QUAD__RCALBG1_CFG4    32'h00000280
`define GTME5_QUAD__RCALBG1_CFG4_SZ 32

`define GTME5_QUAD__RCALBG1_CFG5    32'h00000281
`define GTME5_QUAD__RCALBG1_CFG5_SZ 32

`define GTME5_QUAD__RXRSTDONE_DIST_SEL    32'h00000282
`define GTME5_QUAD__RXRSTDONE_DIST_SEL_SZ 32

`define GTME5_QUAD__SIM_VERSION    32'h00000283
`define GTME5_QUAD__SIM_VERSION_SZ 3

`define GTME5_QUAD__STAT_NPI_REG_LIST    32'h00000284
`define GTME5_QUAD__STAT_NPI_REG_LIST_SZ 32

`define GTME5_QUAD__TERMPROG_CFG    32'h00000285
`define GTME5_QUAD__TERMPROG_CFG_SZ 32

`define GTME5_QUAD__TXRSTDONE_DIST_SEL    32'h00000286
`define GTME5_QUAD__TXRSTDONE_DIST_SEL_SZ 32

`define GTME5_QUAD__UB_CFG0    32'h00000287
`define GTME5_QUAD__UB_CFG0_SZ 32

`endif  // B_GTME5_QUAD_DEFINES_VH