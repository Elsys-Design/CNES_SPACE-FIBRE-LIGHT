// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP48E5_DEFINES_VH
`else
`define B_DSP48E5_DEFINES_VH

// Look-up table parameters
//

`define DSP48E5_ADDR_N  46
`define DSP48E5_ADDR_SZ 32
`define DSP48E5_DATA_SZ 120

// Attribute addresses
//

`define DSP48E5__ACASCREG    32'h00000000
`define DSP48E5__ACASCREG_SZ 32

`define DSP48E5__ADREG    32'h00000001
`define DSP48E5__ADREG_SZ 32

`define DSP48E5__ALUMODEREG    32'h00000002
`define DSP48E5__ALUMODEREG_SZ 32

`define DSP48E5__AMULTSEL    32'h00000003
`define DSP48E5__AMULTSEL_SZ 16

`define DSP48E5__AREG    32'h00000004
`define DSP48E5__AREG_SZ 32

`define DSP48E5__AUTORESET_PATDET    32'h00000005
`define DSP48E5__AUTORESET_PATDET_SZ 120

`define DSP48E5__AUTORESET_PRIORITY    32'h00000006
`define DSP48E5__AUTORESET_PRIORITY_SZ 40

`define DSP48E5__A_INPUT    32'h00000007
`define DSP48E5__A_INPUT_SZ 56

`define DSP48E5__BCASCREG    32'h00000008
`define DSP48E5__BCASCREG_SZ 32

`define DSP48E5__BMULTSEL    32'h00000009
`define DSP48E5__BMULTSEL_SZ 16

`define DSP48E5__BREG    32'h0000000a
`define DSP48E5__BREG_SZ 32

`define DSP48E5__B_INPUT    32'h0000000b
`define DSP48E5__B_INPUT_SZ 56

`define DSP48E5__CARRYINREG    32'h0000000c
`define DSP48E5__CARRYINREG_SZ 32

`define DSP48E5__CARRYINSELREG    32'h0000000d
`define DSP48E5__CARRYINSELREG_SZ 32

`define DSP48E5__CREG    32'h0000000e
`define DSP48E5__CREG_SZ 32

`define DSP48E5__DREG    32'h0000000f
`define DSP48E5__DREG_SZ 32

`define DSP48E5__INMODEREG    32'h00000010
`define DSP48E5__INMODEREG_SZ 32

`define DSP48E5__IS_ALUMODE_INVERTED    32'h00000011
`define DSP48E5__IS_ALUMODE_INVERTED_SZ 4

`define DSP48E5__IS_CARRYIN_INVERTED    32'h00000012
`define DSP48E5__IS_CARRYIN_INVERTED_SZ 1

`define DSP48E5__IS_CLK_INVERTED    32'h00000013
`define DSP48E5__IS_CLK_INVERTED_SZ 1

`define DSP48E5__IS_INMODE_INVERTED    32'h00000014
`define DSP48E5__IS_INMODE_INVERTED_SZ 5

`define DSP48E5__IS_OPMODE_INVERTED    32'h00000015
`define DSP48E5__IS_OPMODE_INVERTED_SZ 9

`define DSP48E5__IS_RSTALLCARRYIN_INVERTED    32'h00000016
`define DSP48E5__IS_RSTALLCARRYIN_INVERTED_SZ 1

`define DSP48E5__IS_RSTALUMODE_INVERTED    32'h00000017
`define DSP48E5__IS_RSTALUMODE_INVERTED_SZ 1

`define DSP48E5__IS_RSTA_INVERTED    32'h00000018
`define DSP48E5__IS_RSTA_INVERTED_SZ 1

`define DSP48E5__IS_RSTB_INVERTED    32'h00000019
`define DSP48E5__IS_RSTB_INVERTED_SZ 1

`define DSP48E5__IS_RSTCTRL_INVERTED    32'h0000001a
`define DSP48E5__IS_RSTCTRL_INVERTED_SZ 1

`define DSP48E5__IS_RSTC_INVERTED    32'h0000001b
`define DSP48E5__IS_RSTC_INVERTED_SZ 1

`define DSP48E5__IS_RSTD_INVERTED    32'h0000001c
`define DSP48E5__IS_RSTD_INVERTED_SZ 1

`define DSP48E5__IS_RSTINMODE_INVERTED    32'h0000001d
`define DSP48E5__IS_RSTINMODE_INVERTED_SZ 1

`define DSP48E5__IS_RSTM_INVERTED    32'h0000001e
`define DSP48E5__IS_RSTM_INVERTED_SZ 1

`define DSP48E5__IS_RSTP_INVERTED    32'h0000001f
`define DSP48E5__IS_RSTP_INVERTED_SZ 1

`define DSP48E5__MASK    32'h00000020
`define DSP48E5__MASK_SZ 48

`define DSP48E5__MREG    32'h00000021
`define DSP48E5__MREG_SZ 32

`define DSP48E5__OPMODEREG    32'h00000022
`define DSP48E5__OPMODEREG_SZ 32

`define DSP48E5__PATTERN    32'h00000023
`define DSP48E5__PATTERN_SZ 48

`define DSP48E5__PREADDINSEL    32'h00000024
`define DSP48E5__PREADDINSEL_SZ 8

`define DSP48E5__PREG    32'h00000025
`define DSP48E5__PREG_SZ 32

`define DSP48E5__RND    32'h00000026
`define DSP48E5__RND_SZ 48

`define DSP48E5__SEL_MASK    32'h00000027
`define DSP48E5__SEL_MASK_SZ 112

`define DSP48E5__SEL_PATTERN    32'h00000028
`define DSP48E5__SEL_PATTERN_SZ 56

`define DSP48E5__USE_MULT    32'h00000029
`define DSP48E5__USE_MULT_SZ 64

`define DSP48E5__USE_PATTERN_DETECT    32'h0000002a
`define DSP48E5__USE_PATTERN_DETECT_SZ 72

`define DSP48E5__USE_SIMD    32'h0000002b
`define DSP48E5__USE_SIMD_SZ 48

`define DSP48E5__USE_WIDEXOR    32'h0000002c
`define DSP48E5__USE_WIDEXOR_SZ 40

`define DSP48E5__XORSIMD    32'h0000002d
`define DSP48E5__XORSIMD_SZ 88

`endif  // B_DSP48E5_DEFINES_VH