-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 02/07/2025
--
-- Description : This is the testbench of the ppl_64_skip_insertion module
----------------------------------------------------------------------------
LIBRARY ieee ;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library work;
use work.pkg_simu.all;

entity tb_ppl_64_skip_insertion is
end entity;

architecture sim of tb_ppl_64_skip_insertion is

  ---------------------------------------------------------
  -----               Component declaration           -----
  ---------------------------------------------------------
  component ppl_64_skip_insertion
   port (
      RST_N                   : in  std_logic;                                          --! global reset
      CLK                     : in  std_logic;                                          --! Clock generated by GTY IP
      -- ppl_64_lane_ctrl_word_insert (PLCWI) Interface
      NEW_DATA_PLCWI          : in  std_logic;                                          --! New data Flag
      DATA_TX_PLCWI           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_PLCWI    : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character from DATA-LINK layer
      WAIT_SEND_DATA_PLSI      : out std_logic;                                          --! Flag to indicates that the lane_ctrl_word_insert send a SKIP control word
      -- HSSL Interface
      DATA_TX_PLSI             : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_PLSI      : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character
      -- ppl_64_lane_init_fsm
      ENABLE_TRANSM_DATA_PLIF : in  std_logic                                           --! Flag to enable to send data
   );
  end component;

  ---------------------------------------------------------
  -----                  Signal declaration           -----
  ---------------------------------------------------------
  -- Inout component
  signal RST_N                   : std_logic := '0';
  signal CLK                     : std_logic := '0';

  signal NEW_DATA_PLCWI          : std_logic                                          := '0';
  signal DATA_TX_PLCWI           : std_logic_vector(C_DATA_LENGTH-1 downto 0)         := (others => '0');
  signal VALID_K_CHARAC_PLCWI    : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0) := (others => '0');
  signal WAIT_SEND_DATA_PLSI      : std_logic;

  signal DATA_TX_PLSI             : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal VALID_K_CHARAC_PLSI      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);

  signal ENABLE_TRANSM_DATA_PLIF : std_logic:='0';
  -- simulation signals
  signal data_2      : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_1      : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_0      : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_2_r    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_1_r    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_0_r    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_2_rr   : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_1_rr   : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');
  signal data_0_rr   : std_logic_vector(C_DATA_LENGTH/2-1 downto 0)        := (others => '0');

  signal k_char_2    : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_1    : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_0    : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_2_r  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_1_r  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_0_r  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_2_rr : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_1_rr : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');
  signal k_char_0_rr : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0):= (others => '0');

  -- Clock generation
  constant CLK_PERIOD : time := 13.334 ns;
  
begin

  ---------------------------------------------------------
  -----                  Instantiation                -----
  ---------------------------------------------------------
  uut: ppl_64_skip_insertion
    port map (
      RST_N                   => RST_N,
      CLK                     => CLK,
      -- ppl_64_lane_ctrl_word_insert (PLCWI) Interface
      NEW_DATA_PLCWI          => NEW_DATA_PLCWI,
      DATA_TX_PLCWI           => DATA_TX_PLCWI,
      VALID_K_CHARAC_PLCWI    => VALID_K_CHARAC_PLCWI,
      WAIT_SEND_DATA_PLSI      => WAIT_SEND_DATA_PLSI,
      -- HSSL Interface
      DATA_TX_PLSI             => DATA_TX_PLSI,
      VALID_K_CHARAC_PLSI      => VALID_K_CHARAC_PLSI,
      -- ppl_64_lane_init_fsm
      ENABLE_TRANSM_DATA_PLIF => ENABLE_TRANSM_DATA_PLIF
    );
  ---------------------------------------------------------
  -----                     Process                   -----
  ---------------------------------------------------------
  clk_process: process
  begin
    while true loop
      CLK <= '0';
      wait for CLK_PERIOD / 2;
      CLK <= '1';
      wait for CLK_PERIOD / 2;
    end loop;
  end process;

  p_reg :process(clk)
  begin
    if rising_edge(clk) then
      data_0      <= data_2;
      k_char_0   <=  k_char_2;

      data_2_r    <= data_2;
      data_2_rr   <= data_2_r;

      data_1_r    <= data_1;
      data_1_rr   <= data_1_r;

      data_0_r    <= data_0;
      data_0_rr   <= data_0_r;

      k_char_2_r  <= k_char_2;
      k_char_2_rr <= k_char_2_r;

      k_char_1_r  <= k_char_1;
      k_char_1_rr <= k_char_1_r;

      k_char_0_r  <= k_char_0;
      k_char_0_rr <= k_char_0_r;
    end if;
  end process p_reg;

  -- Stimulus process
  stim_proc: process
    variable test_failed : boolean := false;
  begin
    -- Reset
    RST_N <= '0';
    wait for 20 ns;
    RST_N <= '1';
    ------------------------------------------------------------
    --                     TX_INIT_ST                         --
    ------------------------------------------------------------
    check_equal("TX_INIT_ST: DATA_TX_PLSI"       , x"0000000000000000", DATA_TX_PLSI,        test_failed);
    check_equal("TX_INIT_ST: VALID_K_CHARAC_PLSI", x"00",               VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_INIT_ST: WAIT_SEND_DATA_PLSI", '0',                 WAIT_SEND_DATA_PLSI, test_failed);
    ------------------------------------------------------------
    --                     TX_DATA_1_ST                       --
    ------------------------------------------------------------
    ENABLE_TRANSM_DATA_PLIF <= '1';
    -- 1st data & k_char generation
    data_1               <= std_logic_vector(to_unsigned(3,C_DATA_LENGTH/2));
    data_2               <= std_logic_vector(to_unsigned(5,C_DATA_LENGTH/2));
    k_char_1             <= std_logic_vector(to_unsigned(1,C_BYTE_BY_WORD_LENGTH/2));
    k_char_2             <= std_logic_vector(to_unsigned(3,C_BYTE_BY_WORD_LENGTH/2));
    DATA_TX_PLCWI        <= data_2 & data_1;
    VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
    wait until rising_edge(clk);
    --2nd data & k_char generation
    data_1               <= std_logic_vector(to_unsigned(6,C_DATA_LENGTH/2));
    data_2               <= std_logic_vector(to_unsigned(10,C_DATA_LENGTH/2));
    k_char_1             <= std_logic_vector(to_unsigned(2,C_BYTE_BY_WORD_LENGTH/2));
    k_char_2             <= std_logic_vector(to_unsigned(6,C_BYTE_BY_WORD_LENGTH/2));
    DATA_TX_PLCWI        <= data_2 & data_1;
    VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
    wait until rising_edge(clk);
    for i in 2 to 2499 loop
      -- data and k_char generation
      data_1               <= std_logic_vector(to_unsigned(i+3,C_DATA_LENGTH/2));
      data_2               <= std_logic_vector(to_unsigned(i+5,C_DATA_LENGTH/2));
      k_char_1             <= std_logic_vector(to_unsigned(i+1,C_BYTE_BY_WORD_LENGTH/2));
      k_char_2             <= std_logic_vector(to_unsigned(i+3,C_BYTE_BY_WORD_LENGTH/2));
      DATA_TX_PLCWI        <= data_2 & data_1;
      VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
      wait until rising_edge(clk);
      -- check outputs
      check_equal("TX_DATA_1_ST: DATA_TX_PLSI i=" & integer'image(i)      , data_2_rr & data_1_rr,     DATA_TX_PLSI,        test_failed);
      check_equal("TX_DATA_1_ST: VALID_K_CHARAC_PLSI i="& integer'image(i), k_char_2_rr & k_char_1_rr, VALID_K_CHARAC_PLSI, test_failed);
      check      ("TX_DATA_1_ST: WAIT_SEND_DATA_PLSI i="& integer'image(i), '0',                       WAIT_SEND_DATA_PLSI, test_failed);
    end loop;
    -- transition state
    -- 1st data & k_char generation for the next 5000 words
    data_1               <= std_logic_vector(to_unsigned(3,C_DATA_LENGTH/2));
    data_2               <= std_logic_vector(to_unsigned(5,C_DATA_LENGTH/2));
    k_char_1             <= std_logic_vector(to_unsigned(1,C_BYTE_BY_WORD_LENGTH/2));
    k_char_2             <= std_logic_vector(to_unsigned(3,C_BYTE_BY_WORD_LENGTH/2));
    DATA_TX_PLCWI        <= data_2 & data_1;
    VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
    wait until rising_edge(clk);
    -- check outputs
    check_equal("TX_DATA_1_ST: DATA_TX_PLSI i=4098",         data_2_rr & data_1_rr,     DATA_TX_PLSI,        test_failed);
    check_equal("TX_DATA_1_ST: VALID_K_CHARAC_PLSI i= 4098", k_char_2_rr & k_char_1_rr, VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_DATA_1_ST: WAIT_SEND_DATA_PLSI i= 4098", '0',                       WAIT_SEND_DATA_PLSI, test_failed);
    --2nd data & k_char generation for the next 5000 words
    data_1               <= std_logic_vector(to_unsigned(6,C_DATA_LENGTH/2));
    data_2               <= std_logic_vector(to_unsigned(10,C_DATA_LENGTH/2));
    k_char_1             <= std_logic_vector(to_unsigned(2,C_BYTE_BY_WORD_LENGTH/2));
    k_char_2             <= std_logic_vector(to_unsigned(6,C_BYTE_BY_WORD_LENGTH/2));
    DATA_TX_PLCWI        <= data_2 & data_1;
    VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
    wait until rising_edge(clk);
    -- check outputs
    check_equal("TX_DATA_1_ST: DATA_TX_PLSI i=4099",         data_2_rr & data_1_rr,     DATA_TX_PLSI,        test_failed);
    check_equal("TX_DATA_1_ST: VALID_K_CHARAC_PLSI i= 4099", k_char_2_rr & k_char_1_rr, VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_DATA_1_ST: WAIT_SEND_DATA_PLSI i= 4099", '0',                       WAIT_SEND_DATA_PLSI, test_failed);
    ------------------------------------------------------------
    --                     TX_SKIP_1_ST                       --
    ------------------------------------------------------------
    --2nd data & k_char generation for the next 5000 words
    data_1               <= std_logic_vector(to_unsigned(9,C_DATA_LENGTH/2));
    data_2               <= std_logic_vector(to_unsigned(15,C_DATA_LENGTH/2));
    k_char_1             <= std_logic_vector(to_unsigned(3,C_BYTE_BY_WORD_LENGTH/2));
    k_char_2             <= std_logic_vector(to_unsigned(9,C_BYTE_BY_WORD_LENGTH/2));
    DATA_TX_PLCWI        <= data_2 & data_1;
    VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
    wait until rising_edge(clk);
    -- check Skip insertion
    check_equal("TX_SKIP_1_ST: DATA_TX_PLSI"       , data_1_rr & C_SKIP_WORD, DATA_TX_PLSI,        test_failed);
    check_equal("TX_SKIP_1_ST: VALID_K_CHARAC_PLSI", k_char_1_rr & x"1",      VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_SKIP_1_ST: WAIT_SEND_DATA_PLSI", '0',                     WAIT_SEND_DATA_PLSI, test_failed);
    ------------------------------------------------------------
    --                     TX_DATA_2_ST                       --
    ------------------------------------------------------------
    for i in 3 to 2500 loop
      -- data and k_char generation
      data_1               <= std_logic_vector(to_unsigned(i+3,C_DATA_LENGTH/2));
      data_2               <= std_logic_vector(to_unsigned(i+5,C_DATA_LENGTH/2));
      k_char_1             <= std_logic_vector(to_unsigned(i+1,C_BYTE_BY_WORD_LENGTH/2));
      k_char_2             <= std_logic_vector(to_unsigned(i+3,C_BYTE_BY_WORD_LENGTH/2));
      DATA_TX_PLCWI        <= data_2 & data_1;
      VALID_K_CHARAC_PLCWI <= k_char_2 & k_char_1;
      wait until rising_edge(clk);
      -- check outputs
      check_equal("TX_DATA_2_ST: DATA_TX_PLSI i=" & integer'image(i)       , data_1_rr & data_0_rr ,    DATA_TX_PLSI,        test_failed);
      check_equal("TX_DATA_2_ST: VALID_K_CHARAC_PLSI i=" & integer'image(i), k_char_1_rr & k_char_0_rr, VALID_K_CHARAC_PLSI, test_failed);
      check      ("TX_DATA_2_ST: WAIT_SEND_DATA_PLSI i=" & integer'image(i), '0',                       WAIT_SEND_DATA_PLSI, test_failed);
    end loop;
    wait until rising_edge(clk);
    -- check outputs and wait send data at '1'
    check_equal("TX_DATA_2_ST: DATA_TX_PLSI i=2500",         data_1_rr & data_0_rr,     DATA_TX_PLSI,        test_failed);
    check_equal("TX_DATA_2_ST: VALID_K_CHARAC_PLSI i= 2500", k_char_1_rr & k_char_0_rr, VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_DATA_2_ST: WAIT_SEND_DATA_PLSI i= 2500", '1',                       WAIT_SEND_DATA_PLSI, test_failed);
    wait until rising_edge(clk);
    ------------------------------------------------------------
    --                     TX_SKIP_2_ST                       --
    ------------------------------------------------------------
    check_equal("TX_SKIP_2_ST: DATA_TX_PLSI"       , C_SKIP_WORD & data_0_rr, DATA_TX_PLSI,        test_failed);
    check_equal("TX_SKIP_2_ST: VALID_K_CHARAC_PLSI", x"1" & k_char_0_rr,      VALID_K_CHARAC_PLSI, test_failed);
    check      ("TX_SKIP_2_ST: WAIT_SEND_DATA_PLSI", '0',                     WAIT_SEND_DATA_PLSI, test_failed);



    log_test_result(test_failed);
    wait;
  end process;

end architecture sim;
