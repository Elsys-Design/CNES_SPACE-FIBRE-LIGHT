// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_ILKNF_DEFINES_VH
`else
`define B_ILKNF_DEFINES_VH

// Look-up table parameters
//

`define ILKNF_ADDR_N  103
`define ILKNF_ADDR_SZ 32
`define ILKNF_DATA_SZ 208

// Attribute addresses
//

`define ILKNF__AXIS_WIDTH    32'h00000000
`define ILKNF__AXIS_WIDTH_SZ 12

`define ILKNF__C0_CTL_RX_AXIS_WIDTH    32'h00000001
`define ILKNF__C0_CTL_RX_AXIS_WIDTH_SZ 3

`define ILKNF__C0_CTL_RX_BURSTMAX    32'h00000002
`define ILKNF__C0_CTL_RX_BURSTMAX_SZ 2

`define ILKNF__C0_CTL_RX_CHAN_EXT    32'h00000003
`define ILKNF__C0_CTL_RX_CHAN_EXT_SZ 2

`define ILKNF__C0_CTL_RX_FECFRAMELEN_MINUS1    32'h00000004
`define ILKNF__C0_CTL_RX_FECFRAMELEN_MINUS1_SZ 12

`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID0    32'h00000005
`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID0_SZ 64

`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID4    32'h00000006
`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID4_SZ 64

`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID5    32'h00000007
`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID5_SZ 64

`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID6    32'h00000008
`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID6_SZ 64

`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID7    32'h00000009
`define ILKNF__C0_CTL_RX_FEC_VL_MARKER_ID7_SZ 64

`define ILKNF__C0_CTL_RX_GEARBOX_MODE    32'h0000000a
`define ILKNF__C0_CTL_RX_GEARBOX_MODE_SZ 2

`define ILKNF__C0_CTL_RX_LAST_LANE    32'h0000000b
`define ILKNF__C0_CTL_RX_LAST_LANE_SZ 5

`define ILKNF__C0_CTL_RX_MFRAMELEN_MINUS1    32'h0000000c
`define ILKNF__C0_CTL_RX_MFRAMELEN_MINUS1_SZ 16

`define ILKNF__C0_CTL_RX_PACKET_MODE    32'h0000000d
`define ILKNF__C0_CTL_RX_PACKET_MODE_SZ 40

`define ILKNF__C0_CTL_RX_RATE_ADAPT_DEC    32'h0000000e
`define ILKNF__C0_CTL_RX_RATE_ADAPT_DEC_SZ 8

`define ILKNF__C0_CTL_RX_RATE_ADAPT_INC    32'h0000000f
`define ILKNF__C0_CTL_RX_RATE_ADAPT_INC_SZ 8

`define ILKNF__C0_CTL_RX_SERDES_INTF_MODE    32'h00000010
`define ILKNF__C0_CTL_RX_SERDES_INTF_MODE_SZ 2

`define ILKNF__C0_CTL_TX_AXIS_WIDTH    32'h00000011
`define ILKNF__C0_CTL_TX_AXIS_WIDTH_SZ 3

`define ILKNF__C0_CTL_TX_BURSTMAX    32'h00000012
`define ILKNF__C0_CTL_TX_BURSTMAX_SZ 2

`define ILKNF__C0_CTL_TX_BURSTSHORT    32'h00000013
`define ILKNF__C0_CTL_TX_BURSTSHORT_SZ 3

`define ILKNF__C0_CTL_TX_CHAN_EXT    32'h00000014
`define ILKNF__C0_CTL_TX_CHAN_EXT_SZ 2

`define ILKNF__C0_CTL_TX_DISABLE_SKIPWORD    32'h00000015
`define ILKNF__C0_CTL_TX_DISABLE_SKIPWORD_SZ 40

`define ILKNF__C0_CTL_TX_FC_CALLEN    32'h00000016
`define ILKNF__C0_CTL_TX_FC_CALLEN_SZ 4

`define ILKNF__C0_CTL_TX_FECFRAMELEN_MINUS1    32'h00000017
`define ILKNF__C0_CTL_TX_FECFRAMELEN_MINUS1_SZ 12

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID0    32'h00000018
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID0_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID1    32'h00000019
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID1_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID10    32'h0000001a
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID10_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID11    32'h0000001b
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID11_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID12    32'h0000001c
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID12_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID13    32'h0000001d
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID13_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID14    32'h0000001e
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID14_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID15    32'h0000001f
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID15_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID16    32'h00000020
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID16_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID17    32'h00000021
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID17_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID18    32'h00000022
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID18_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID19    32'h00000023
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID19_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID2    32'h00000024
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID2_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID3    32'h00000025
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID3_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID4    32'h00000026
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID4_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID5    32'h00000027
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID5_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID6    32'h00000028
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID6_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID7    32'h00000029
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID7_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID8    32'h0000002a
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID8_SZ 64

`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID9    32'h0000002b
`define ILKNF__C0_CTL_TX_FEC_VL_MARKER_ID9_SZ 64

`define ILKNF__C0_CTL_TX_GEARBOX_MODE    32'h0000002c
`define ILKNF__C0_CTL_TX_GEARBOX_MODE_SZ 2

`define ILKNF__C0_CTL_TX_LAST_LANE    32'h0000002d
`define ILKNF__C0_CTL_TX_LAST_LANE_SZ 5

`define ILKNF__C0_CTL_TX_MFRAMELEN_MINUS1    32'h0000002e
`define ILKNF__C0_CTL_TX_MFRAMELEN_MINUS1_SZ 16

`define ILKNF__C0_CTL_TX_RDYOUT_THRESH    32'h0000002f
`define ILKNF__C0_CTL_TX_RDYOUT_THRESH_SZ 4

`define ILKNF__C0_CTL_TX_RLIM_DELTA    32'h00000030
`define ILKNF__C0_CTL_TX_RLIM_DELTA_SZ 16

`define ILKNF__C0_CTL_TX_RLIM_ENABLE    32'h00000031
`define ILKNF__C0_CTL_TX_RLIM_ENABLE_SZ 40

`define ILKNF__C0_CTL_TX_RLIM_MAX    32'h00000032
`define ILKNF__C0_CTL_TX_RLIM_MAX_SZ 16

`define ILKNF__C0_CTL_TX_SERDES_INTF_MODE    32'h00000033
`define ILKNF__C0_CTL_TX_SERDES_INTF_MODE_SZ 2

`define ILKNF__CORE_MODE    32'h00000034
`define ILKNF__CORE_MODE_SZ 120

`define ILKNF__CTL_CORE_MODE    32'h00000035
`define ILKNF__CTL_CORE_MODE_SZ 2

`define ILKNF__CTL_REVISION    32'h00000036
`define ILKNF__CTL_REVISION_SZ 32

`define ILKNF__CTL_RSVD2_IN    32'h00000037
`define ILKNF__CTL_RSVD2_IN_SZ 32

`define ILKNF__CTL_RX_AXI_SHUTDOWN_GATE    32'h00000038
`define ILKNF__CTL_RX_AXI_SHUTDOWN_GATE_SZ 1

`define ILKNF__CTL_RX_CORE_SHUTDOWN_GATE    32'h00000039
`define ILKNF__CTL_RX_CORE_SHUTDOWN_GATE_SZ 1

`define ILKNF__CTL_RX_DEBUG_SELECT    32'h0000003a
`define ILKNF__CTL_RX_DEBUG_SELECT_SZ 6

`define ILKNF__CTL_RX_FEC0_SLICE0_MODE    32'h0000003b
`define ILKNF__CTL_RX_FEC0_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC0_SLICE1_MODE    32'h0000003c
`define ILKNF__CTL_RX_FEC0_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC1_SLICE0_MODE    32'h0000003d
`define ILKNF__CTL_RX_FEC1_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC1_SLICE1_MODE    32'h0000003e
`define ILKNF__CTL_RX_FEC1_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC2_SLICE0_MODE    32'h0000003f
`define ILKNF__CTL_RX_FEC2_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC2_SLICE1_MODE    32'h00000040
`define ILKNF__CTL_RX_FEC2_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC3_SLICE0_MODE    32'h00000041
`define ILKNF__CTL_RX_FEC3_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC3_SLICE1_MODE    32'h00000042
`define ILKNF__CTL_RX_FEC3_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC4_SLICE0_MODE    32'h00000043
`define ILKNF__CTL_RX_FEC4_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC4_SLICE1_MODE    32'h00000044
`define ILKNF__CTL_RX_FEC4_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC5_SLICE0_MODE    32'h00000045
`define ILKNF__CTL_RX_FEC5_SLICE0_MODE_SZ 2

`define ILKNF__CTL_RX_FEC5_SLICE1_MODE    32'h00000046
`define ILKNF__CTL_RX_FEC5_SLICE1_MODE_SZ 2

`define ILKNF__CTL_RX_FEC_ONLY_ENABLE    32'h00000047
`define ILKNF__CTL_RX_FEC_ONLY_ENABLE_SZ 2

`define ILKNF__CTL_RX_LANE_SHUTDOWN_GATE    32'h00000048
`define ILKNF__CTL_RX_LANE_SHUTDOWN_GATE_SZ 6

`define ILKNF__CTL_TX_AXI_SHUTDOWN_GATE    32'h00000049
`define ILKNF__CTL_TX_AXI_SHUTDOWN_GATE_SZ 1

`define ILKNF__CTL_TX_CORE_SHUTDOWN_GATE    32'h0000004a
`define ILKNF__CTL_TX_CORE_SHUTDOWN_GATE_SZ 1

`define ILKNF__CTL_TX_DEBUG_SELECT    32'h0000004b
`define ILKNF__CTL_TX_DEBUG_SELECT_SZ 6

`define ILKNF__CTL_TX_FEC0_SLICE0_MODE    32'h0000004c
`define ILKNF__CTL_TX_FEC0_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC0_SLICE1_MODE    32'h0000004d
`define ILKNF__CTL_TX_FEC0_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC1_SLICE0_MODE    32'h0000004e
`define ILKNF__CTL_TX_FEC1_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC1_SLICE1_MODE    32'h0000004f
`define ILKNF__CTL_TX_FEC1_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC2_SLICE0_MODE    32'h00000050
`define ILKNF__CTL_TX_FEC2_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC2_SLICE1_MODE    32'h00000051
`define ILKNF__CTL_TX_FEC2_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC3_SLICE0_MODE    32'h00000052
`define ILKNF__CTL_TX_FEC3_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC3_SLICE1_MODE    32'h00000053
`define ILKNF__CTL_TX_FEC3_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC4_SLICE0_MODE    32'h00000054
`define ILKNF__CTL_TX_FEC4_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC4_SLICE1_MODE    32'h00000055
`define ILKNF__CTL_TX_FEC4_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC5_SLICE0_MODE    32'h00000056
`define ILKNF__CTL_TX_FEC5_SLICE0_MODE_SZ 2

`define ILKNF__CTL_TX_FEC5_SLICE1_MODE    32'h00000057
`define ILKNF__CTL_TX_FEC5_SLICE1_MODE_SZ 2

`define ILKNF__CTL_TX_FEC_ONLY_ENABLE    32'h00000058
`define ILKNF__CTL_TX_FEC_ONLY_ENABLE_SZ 2

`define ILKNF__CTL_TX_LANE_SHUTDOWN_GATE    32'h00000059
`define ILKNF__CTL_TX_LANE_SHUTDOWN_GATE_SZ 6

`define ILKNF__FEC    32'h0000005a
`define ILKNF__FEC_SZ 64

`define ILKNF__FEC_FOR_ILKN_LANES    32'h0000005b
`define ILKNF__FEC_FOR_ILKN_LANES_SZ 96

`define ILKNF__FEC_ONLY_ENABLE    32'h0000005c
`define ILKNF__FEC_ONLY_ENABLE_SZ 160

`define ILKNF__FEC_ONLY_MULT_FACTOR    32'h0000005d
`define ILKNF__FEC_ONLY_MULT_FACTOR_SZ 64

`define ILKNF__GEARBOX_MODE    32'h0000005e
`define ILKNF__GEARBOX_MODE_SZ 80

`define ILKNF__ILKN_LANE_SERIAL_RATE    32'h0000005f
`define ILKNF__ILKN_LANE_SERIAL_RATE_SZ 64

`define ILKNF__ILKN_MODE    32'h00000060
`define ILKNF__ILKN_MODE_SZ 208

`define ILKNF__LANE_CONNECTIVITY    32'h00000061
`define ILKNF__LANE_CONNECTIVITY_SZ 32

`define ILKNF__MEM_CTRL    32'h00000062
`define ILKNF__MEM_CTRL_SZ 8

`define ILKNF__NUM_100G_FEC_NOILKN_PORTS    32'h00000063
`define ILKNF__NUM_100G_FEC_NOILKN_PORTS_SZ 3

`define ILKNF__NUM_50G_FEC_NOILKN_PORTS    32'h00000064
`define ILKNF__NUM_50G_FEC_NOILKN_PORTS_SZ 4

`define ILKNF__NUM_ILKN_SERDES_LANES    32'h00000065
`define ILKNF__NUM_ILKN_SERDES_LANES_SZ 5

`define ILKNF__SIM_VERSION    32'h00000066
`define ILKNF__SIM_VERSION_SZ 4

`endif  // B_ILKNF_DEFINES_VH