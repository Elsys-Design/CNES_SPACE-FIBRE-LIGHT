// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_X5PLL_DEFINES_VH
`else
`define B_X5PLL_DEFINES_VH

// Look-up table parameters
//

`define X5PLL_ADDR_N  52
`define X5PLL_ADDR_SZ 32
`define X5PLL_DATA_SZ 64

// Attribute addresses
//

`define X5PLL__CLKFBOUT_MULT    32'h00000000
`define X5PLL__CLKFBOUT_MULT_SZ 32

`define X5PLL__CLKFBOUT_PHASE    32'h00000001
`define X5PLL__CLKFBOUT_PHASE_SZ 64

`define X5PLL__CLKIN_FREQ_MAX    32'h00000002
`define X5PLL__CLKIN_FREQ_MAX_SZ 64

`define X5PLL__CLKIN_FREQ_MIN    32'h00000003
`define X5PLL__CLKIN_FREQ_MIN_SZ 64

`define X5PLL__CLKIN_PERIOD    32'h00000004
`define X5PLL__CLKIN_PERIOD_SZ 64

`define X5PLL__CLKOUT0_DIVIDE    32'h00000005
`define X5PLL__CLKOUT0_DIVIDE_SZ 32

`define X5PLL__CLKOUT0_DUTY_CYCLE    32'h00000006
`define X5PLL__CLKOUT0_DUTY_CYCLE_SZ 64

`define X5PLL__CLKOUT0_PHASE    32'h00000007
`define X5PLL__CLKOUT0_PHASE_SZ 64

`define X5PLL__CLKOUT0_PHASE_CTRL    32'h00000008
`define X5PLL__CLKOUT0_PHASE_CTRL_SZ 2

`define X5PLL__CLKOUT1_DIVIDE    32'h00000009
`define X5PLL__CLKOUT1_DIVIDE_SZ 32

`define X5PLL__CLKOUT1_DUTY_CYCLE    32'h0000000a
`define X5PLL__CLKOUT1_DUTY_CYCLE_SZ 64

`define X5PLL__CLKOUT1_PHASE    32'h0000000b
`define X5PLL__CLKOUT1_PHASE_SZ 64

`define X5PLL__CLKOUT1_PHASE_CTRL    32'h0000000c
`define X5PLL__CLKOUT1_PHASE_CTRL_SZ 2

`define X5PLL__CLKOUT2_DIVIDE    32'h0000000d
`define X5PLL__CLKOUT2_DIVIDE_SZ 32

`define X5PLL__CLKOUT2_DUTY_CYCLE    32'h0000000e
`define X5PLL__CLKOUT2_DUTY_CYCLE_SZ 64

`define X5PLL__CLKOUT2_PHASE    32'h0000000f
`define X5PLL__CLKOUT2_PHASE_SZ 64

`define X5PLL__CLKOUT2_PHASE_CTRL    32'h00000010
`define X5PLL__CLKOUT2_PHASE_CTRL_SZ 2

`define X5PLL__CLKOUT3_DIVIDE    32'h00000011
`define X5PLL__CLKOUT3_DIVIDE_SZ 32

`define X5PLL__CLKOUT3_DUTY_CYCLE    32'h00000012
`define X5PLL__CLKOUT3_DUTY_CYCLE_SZ 64

`define X5PLL__CLKOUT3_PHASE    32'h00000013
`define X5PLL__CLKOUT3_PHASE_SZ 64

`define X5PLL__CLKOUT3_PHASE_CTRL    32'h00000014
`define X5PLL__CLKOUT3_PHASE_CTRL_SZ 2

`define X5PLL__CLKOUTPHY_CASCIN_EN    32'h00000015
`define X5PLL__CLKOUTPHY_CASCIN_EN_SZ 1

`define X5PLL__CLKOUTPHY_CASCOUT_EN    32'h00000016
`define X5PLL__CLKOUTPHY_CASCOUT_EN_SZ 1

`define X5PLL__CLKOUTPHY_DIVIDE    32'h00000017
`define X5PLL__CLKOUTPHY_DIVIDE_SZ 40

`define X5PLL__CLKPFD_FREQ_MAX    32'h00000018
`define X5PLL__CLKPFD_FREQ_MAX_SZ 64

`define X5PLL__CLKPFD_FREQ_MIN    32'h00000019
`define X5PLL__CLKPFD_FREQ_MIN_SZ 64

`define X5PLL__DESKEW2_MUXIN_SEL    32'h0000001a
`define X5PLL__DESKEW2_MUXIN_SEL_SZ 1

`define X5PLL__DESKEW_DELAY1    32'h0000001b
`define X5PLL__DESKEW_DELAY1_SZ 32

`define X5PLL__DESKEW_DELAY2    32'h0000001c
`define X5PLL__DESKEW_DELAY2_SZ 32

`define X5PLL__DESKEW_DELAY_EN1    32'h0000001d
`define X5PLL__DESKEW_DELAY_EN1_SZ 40

`define X5PLL__DESKEW_DELAY_EN2    32'h0000001e
`define X5PLL__DESKEW_DELAY_EN2_SZ 40

`define X5PLL__DESKEW_DELAY_PATH1    32'h0000001f
`define X5PLL__DESKEW_DELAY_PATH1_SZ 40

`define X5PLL__DESKEW_DELAY_PATH2    32'h00000020
`define X5PLL__DESKEW_DELAY_PATH2_SZ 40

`define X5PLL__DESKEW_MUXIN_SEL    32'h00000021
`define X5PLL__DESKEW_MUXIN_SEL_SZ 1

`define X5PLL__DIV4_CLKOUT012    32'h00000022
`define X5PLL__DIV4_CLKOUT012_SZ 1

`define X5PLL__DIV4_CLKOUT3    32'h00000023
`define X5PLL__DIV4_CLKOUT3_SZ 1

`define X5PLL__DIVCLK_DIVIDE    32'h00000024
`define X5PLL__DIVCLK_DIVIDE_SZ 32

`define X5PLL__IS_CLKFB1_DESKEW_INVERTED    32'h00000025
`define X5PLL__IS_CLKFB1_DESKEW_INVERTED_SZ 1

`define X5PLL__IS_CLKFB2_DESKEW_INVERTED    32'h00000026
`define X5PLL__IS_CLKFB2_DESKEW_INVERTED_SZ 1

`define X5PLL__IS_CLKIN1_DESKEW_INVERTED    32'h00000027
`define X5PLL__IS_CLKIN1_DESKEW_INVERTED_SZ 1

`define X5PLL__IS_CLKIN2_DESKEW_INVERTED    32'h00000028
`define X5PLL__IS_CLKIN2_DESKEW_INVERTED_SZ 1

`define X5PLL__IS_CLKIN_INVERTED    32'h00000029
`define X5PLL__IS_CLKIN_INVERTED_SZ 1

`define X5PLL__IS_PSEN_INVERTED    32'h0000002a
`define X5PLL__IS_PSEN_INVERTED_SZ 1

`define X5PLL__IS_PSINCDEC_INVERTED    32'h0000002b
`define X5PLL__IS_PSINCDEC_INVERTED_SZ 1

`define X5PLL__IS_PWRDWN_INVERTED    32'h0000002c
`define X5PLL__IS_PWRDWN_INVERTED_SZ 1

`define X5PLL__IS_RST_INVERTED    32'h0000002d
`define X5PLL__IS_RST_INVERTED_SZ 1

`define X5PLL__LOCK_WAIT    32'h0000002e
`define X5PLL__LOCK_WAIT_SZ 40

`define X5PLL__REF_JITTER    32'h0000002f
`define X5PLL__REF_JITTER_SZ 64

`define X5PLL__SIM_ADJ_CLK0_CASCADE    32'h00000030
`define X5PLL__SIM_ADJ_CLK0_CASCADE_SZ 40

`define X5PLL__VCOCLK_FREQ_MAX    32'h00000031
`define X5PLL__VCOCLK_FREQ_MAX_SZ 64

`define X5PLL__VCOCLK_FREQ_MIN    32'h00000032
`define X5PLL__VCOCLK_FREQ_MIN_SZ 64

`define X5PLL__XPLL_CONNECT_TO_NOCMC    32'h00000033
`define X5PLL__XPLL_CONNECT_TO_NOCMC_SZ 32

`endif  // B_X5PLL_DEFINES_VH