-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibre_Light Versal target
--
-- Creation date : 04/08/2025
--
-- Description : This module implement the Physical and Lane layer of an IP
-- SpaceFibre Light.
-- The Physical layer is carried by an NanoXplore IP
-- The Lane layer is carried by owner's code and an NanoXplore IP
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity phy_plus_lane_64b is
  port(
    RST_N                            : in  std_logic;                       --! Global reset. Active Low
    CLK                              : in  std_logic;                       --! Main clock
    -- Reset_gen interface
    LANE_RESET_PPL_OUT               : out std_logic;
    RST_TXCLK_N                      : in  std_logic;                       --! Synchronous reset on clock generated by GTY PLL
    CLK_TX_OUT                       : out std_logic;                       --! Clock generated by manufacturer IP
    RST_TX_DONE                      : out std_logic;                       --! Up when internal rx reset done
    -- CLK HSSL signals
    CLK_REF_N                        : in std_logic;                        --! Referance HSSL IP Clock (neg)
    CLK_REF_P                        : in std_logic;                        --! Referance HSSL IP Clock (pos)
    -- FROM Data-link layer
    DATA_TX                          : in  std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be send from Data-Link Layer
    LANE_RESET_DL                    : in  std_logic;                       --! Lane reset command from Data-Link Layer
    CAPABILITY_TX                    : in  std_logic_vector(07 downto 00);  --! Capability field send in INIT3 control word
    NEW_DATA_TX                      : in  std_logic;                       --! Flag new data
    VALID_K_CHARAC_TX                : in  std_logic_vector(03 downto 00);  --! 4-bit valid K character flags from Data-link layer
    FIFO_TX_FULL                     : out std_logic;                       --! FiFo TX full flag

    -- TO Data-link layer
    FIFO_RX_RD_EN                    : in  std_logic;                       --! FiFo RX read enable flag
    DATA_RX                          : out std_logic_vector(31 downto 00);  --! 32-bit Data parallel to be received to Data-Link Layer
    FIFO_RX_EMPTY                    : out std_logic;                       --! FiFo RX empty flag
    FIFO_RX_DATA_VALID               : out std_logic;                       --! FiFo RX data valid flag
    VALID_K_CHARAC_RX                : out std_logic_vector(03 downto 00);  --! 4-bit valid K character flags to Data-link layer
    FAR_END_CAPA_DL                  : out std_logic_vector(07 downto 00);  --! Capability field receive in INIT3 control word
    LANE_ACTIVE_DL                   : out std_logic;                       --! Lane Active flag for the DATA Link Layer

    -- FROM/TO Outside
    TX_POS                           : out std_logic;                       --! Positive LVDS serial data send
    TX_NEG                           : out std_logic;                       --! Negative LVDS serial data send
    RX_POS                           : in  std_logic;                       --! Positive LVDS serial data received
    RX_NEG                           : in  std_logic;                       --! Negative LVDS serial data received

    -- PARAMETERS and STATUS
    LANE_START                       : in  std_logic;                       --! Asserts or de-asserts LaneStart for the lane
    AUTOSTART                        : in  std_logic;                       --! Asserts or de-asserts AutoStart for the lane
    LANE_RESET                       : in  std_logic;                       --! Asserts or de-asserts LaneReset for the lane
    PARALLEL_LOOPBACK_EN             : in  std_logic;                       --! Enables or disables the parallel loopback for the lane
    STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  --! In case of error, pauses communication
    NEAR_END_SERIAL_LB_EN            : in  std_logic;                       --! Enables or disables the near-end serial loopback for the lane
    FAR_END_SERIAL_LB_EN             : in  std_logic;                       --! Enables or disables the far-end serial loopback for the lane

    LANE_STATE                       : out std_logic_vector(03 downto 00);  --! Indicates the current state of the Lane Initialization state machine in a lane
    RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  --! Counter of error detected on the RX link
    RX_ERROR_OVF                     : out std_logic;                       --! Overflow flag of the RX_ERROR_CNT
    LOSS_SIGNAL                      : out std_logic;                       --! Set when no signal is received on RX link
    FAR_END_CAPA                     : out std_logic_vector(07 downto 00);  --! Capabilities field (INT3 flags)
    RX_POLARITY                      : out std_logic                        --! Set when the receiver polarity is inverted
  );
end phy_plus_lane_64b;

architecture rtl of phy_plus_lane_64b is
---------------------------------------------------------
-----               Component declaration           -----
---------------------------------------------------------
-- HSSL
  component SpaceFibre_64b
    port (
      HSSL_CLOCK_I                  : in  std_logic_vector(3 downto 0);
      RX0N                          : in  std_logic;
      RX0P                          : in  std_logic;
      RX1N                          : in  std_logic;
      RX1P                          : in  std_logic;
      RX2N                          : in  std_logic;
      RX2P                          : in  std_logic;
      RX3N                          : in  std_logic;
      RX3P                          : in  std_logic;
      TX0N                          : out std_logic;
      TX0P                          : out std_logic;
      TX1N                          : out std_logic;
      TX1P                          : out std_logic;
      TX2N                          : out std_logic;
      TX2P                          : out std_logic;
      TX3N                          : out std_logic;
      TX3P                          : out std_logic;
      CKREFN                        : in  std_logic;
      CKREFP                        : in  std_logic;
      CLOCK_O                       : out std_logic;
      DYN_CFG_EN_I                  : in  std_logic;
      DYN_ADDR_I                    : in  std_logic_vector(3 downto 0);
      DYN_CALIBRATION_CS_N_I        : in  std_logic;
      DYN_LANE_CS_N_I               : in  std_logic_vector(3 downto 0);
      DYN_WDATA_I                   : in  std_logic_vector(11 downto 0);
      DYN_WDATA_SEL_I               : in  std_logic;
      DYN_WE_N_I                    : in  std_logic;
      PLL_PMA_LOCK_ANALOG           : out std_logic;
      PLL_PMA_PWR_UP_I              : in  std_logic;
      PLL_PMA_RST_N_I               : in  std_logic;
      PLL_LOCK                      : out std_logic;
      TX0_BUSY_O                    : out std_logic;
      TX0_CLK_ENA_I                 : in  std_logic;
      TX0_CLK_O                     : out std_logic;
      TX0_DATA_I                    : in  std_logic_vector(63 downto 0);
      TX0_CTRL_DRIVER_PWRDWN_N_I    : in  std_logic;
      TX0_RST_N_I                   : in  std_logic;
      TX0_CTRL_CHAR_IS_K_I          : in  std_logic_vector(7 downto 0);
      RX0_BUSY_O                    : out std_logic;
      RX0_CTRL_EL_BUFF_STAT_O       : out std_logic_vector (7 downto 0);
      RX0_CTRL_CHAR_IS_ALIGNED_O    : out std_logic;
      RX0_CTRL_CHAR_IS_COMMA_O      : out std_logic_vector(7 downto 0);
      RX0_CTRL_CHAR_IS_F_O          : out std_logic_vector(7 downto 0);
      RX0_CTRL_CHAR_IS_K_O          : out std_logic_vector(7 downto 0);
      RX0_CTRL_DISP_ERR_O           : out std_logic_vector(7 downto 0);
      RX0_CTRL_NOT_IN_TABLE_O       : out std_logic_vector(7 downto 0);
      RX0_CTRL_VALID_REALIGN_O      : out std_logic;
      RX0_DATA_O                    : out std_logic_vector(63 downto 0);
      RX0_OVS_BIT_SEL_I             : in  std_logic_vector(1 downto 0);
      RX0_EYE_RST_I                 : in  std_logic;
      RX0_PMA_LL_FAST_LOCKED_O      : out std_logic;
      RX0_PMA_LL_SLOW_LOCKED_O      : out std_logic;
      RX0_PMA_LOSS_OF_SIGNAL_O      : out std_logic;
      RX0_PMA_PLL_LOCK_O            : out std_logic;
      RX0_PMA_PLL_LOCK_TRACK_O      : out std_logic;
      RX0_PMA_RST_N_I               : in  std_logic;
      RX0_PMA_PWR_UP_I              : in  std_logic;
      RX0_RST_N_I                   : in  std_logic;
      RX0_TEST_O                    : out std_logic_vector (7 downto 0);
      RX0_REPLACE_EN_I              : in  std_logic;
      RX0_ALIGN_SYNC_I              : in  std_logic;
      RX0_EL_BUFF_RST_I             : in  std_logic
    );
  end component;

  component ppl_64_init_hssl
    port (
      RST_N                            : in  std_logic; --! Global reset, Active Low
      CLK                              : in  std_logic; --! Clock generated by HSSL IP
      -- ppl_64_lane_init_fsm (PLIF) interface
      RECEIVER_DISABLED_PLIF           : in std_logic;  --! Flag to enable RX function of HSSL IP
      CDR_PLIF                         : in std_logic;  --! Flag to enable CDR_PLIF function of HSSL IP
      TRANSMITTER_DISABLED_PLIF        : in std_logic;  --! Flag to enable TX function of HSSL IP
      -- HSSL interface
      PLL_PMA_PWR_UP_PLIH              : out std_logic; --! '0’- PLL is disabled. Dynamic power consumption is highly reduced. ‘1’ - PLL is active. Normal PLL operation
      TX_DRIVER_PWRDWN_N_PLIH          : out std_logic; --! TX driver is powered down (TX lanes stay at high impedance) , when asserted. Active low
      PLL_PMA_RST_N_PLIH               : out std_logic; --! Active-low PMA PLL reset
      PLL_PMA_LOCK_ANALOG_HSSL         : in  std_logic; --! PMA PLL is locked (Analog Signal)
      TX_RST_N_PLIH                    : out std_logic; --! TX PCS reset. Active low
      TX_BUSY_HSSL                     : in  std_logic; --! Indicates that RX PCS is busy while being reset
      RX_PMA_PWR_UP_PLIH               : out std_logic; --! Resets RX PLL and CDR, when asserted. Active low.
      RX_PMA_RST_N_PLIH                : out std_logic; --! RX PCS reset. Active low
      RX_PMA_LL_SLOW_LOCKED_HSSL       : in  std_logic; --! Asserted when RX PMA Lead Lag (LL) PLL is locked.
      RX_RST_N_PLIH                    : out std_logic; --! PMA PLL power up
      RX_BUSY_HSSL                     : in  std_logic; --! Indicates that RX PCS is busy while being reseted
      -- Output
      HSSL_RESET_DONE_PLIH             : out std_logic  --! HSSL reset done flag
    );
  end component;

  -- TX FLOW
  component ppl_64_bus_concat_tx
    port (
      RST_N                        : in  std_logic;                                   --! global reset
      CLK                          : in  std_logic;                                   --! Clock synchronous with the Data-Link Layer
      -- Data-link layer interface
      DATA_TX_DL                   : in  std_logic_vector(31 downto 0);               --! 32-bit data parallel to be sent from Data-Link Layer
      NEW_DATA_TX_DL               : in  std_logic;                                   --! New data flag
      VALID_K_CHARAC_TX_DL         : in  std_logic_vector(3 downto 0);                --! 4-bit valid K character flags from Data-link layer
      CAPABILITY_TX_DL             : in  std_logic_vector(7 downto 0);                --! Capability field sent in INIT3 control word
      LANE_RESET_DL                : in  std_logic;                                   --! Lane reset command from Data-Link Layer
      -- ppl_64_data_fifo_tx (PLDFT) interface
      DATA_TX_PLBCT                : out std_logic_vector(C_DATA_WIDTH-1  downto 0);  --! 64-bit Data parallel to be sent
      NEW_DATA_TX_PLBCT            : out std_logic;                                   --! New data flag
      VALID_K_CHARAC_TX_PLBCT      : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags
      -- ppl_64_ctrl_fifo_tx (PLCFT) interface
      CAPABILITY_TX_PLBCT          : out std_logic_vector(7 downto 0);                --! Capability field sent in INIT3 control word
      LANE_RESET_PLBCT             : out std_logic                                    --! Lane reset command
    );
  end component;

  component ppl_64_lane_ctrl_word_insert
    port (
      RST_N                                : in  std_logic;                                   --! Global reset Active Low
      CLK                                  : in  std_logic;                                   --! Clock generated by HSSL IP
      -- Data-Link interface
      RD_DATA_EN_PLCWI                     : out std_logic;                                   --! Read command to receive data from the Data-Link layer
      RD_DATA_VALID_DL                     : in  std_logic;                                   --! Data valid flag from the Data-Link layer
      CAPABILITY_DL                        : in  std_logic_vector(7 downto 0);                --! Capability field from the Data-Link layer
      DATA_TX_DL                           : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data received from the Data-Link layer
      VALID_K_CHARAC_DL                    : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicating which bytes are K characters from the Data-Link layer
      NO_DATA_DL                           : in  std_logic;                                   --! Flag enabling IDLE word insertion when no data is available from the Data-Link layer
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI                  : in  std_logic;                                   --! Flag indicating that skip_insertion is sending a SKIP control word
      NEW_DATA_PLCWI                       : out std_logic;                                   --! New data available for skip_insertion
      DATA_TX_PLCWI                        : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to be sent to the physical layer
      VALID_K_CHARAC_PLCWI                 : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicating which bytes are K characters
      -- ppl_64_lane_init_fsm (PLIF) interface
      SEND_INIT1_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT1 control word followed by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT2 control word followed by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD_PLIF            : in  std_logic;                                   --! Flag to send INIT3 control word followed by 64 pseudo-random data words
      ENABLE_TRANSM_DATA_PLIF              : in  std_logic;                                   --! Flag to enable data transmission
      SEND_32_STANDBY_CTRL_WORDS_PLIF      : in  std_logic;                                   --! Flag to send 32 STANDBY control words
      SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF  : in  std_logic;                                   --! Flag to send 32 LOSS_SIGNAL control words
      STANDBY_SIGNAL_X32_PLCWI             : out std_logic;                                   --! Flag indicating 32 STANDBY control words have been sent
      LOST_SIGNAL_X32_PLCWI                : out std_logic;                                   --! Flag indicating 32 LOSS_SIGNAL control words have been sent
      LOST_CAUSE_PLIF                      : in  std_logic_vector(1 downto 0);                --! Indicates the reason for LOST_SIGNAL
      -- MIB interface
      STANDBY_REASON_MIB                   : in  std_logic_vector(7 downto 0)                 --! Standby reason from MIB
    );
  end component;

  component ppl_64_skip_insertion
    port (
      RST_N                   : in  std_logic;                                   --! Global reset (Active low)
      CLK                     : in  std_logic;                                   --! Clock generated by HSSL IP
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      NEW_DATA_PLCWI          : in  std_logic;                                   --! New data Flag
      DATA_TX_PLCWI           : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! Data 64-bit received from DATA_LINK layer
      VALID_K_CHARAC_PLCWI    : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicate which byte is a K character from DATA-LINK layer
      WAIT_SEND_DATA_PLSI     : out std_logic;                                   --! Flag to indicate that the lane_ctrl_word_insert sends a SKIP control word
      -- HSSL interface
      DATA_TX_PLSI            : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! Data 64-bit sent to manufacturer IP
      VALID_K_CHARAC_PLSI     : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flags indicate which byte is a K character
      -- ppl_64_lane_init_fsm (PLIF) interface
      ENABLE_TRANSM_DATA_PLIF : in  std_logic                                    --! Flag to enable sending data
    );
  end component;

  component ppl_64_parallel_loopback
    port (
      CLK                      : in  std_logic;                                   --! Clock generated by HSSL IP
      RST_N                    : in  std_logic;                                   --! Global reset. Active low
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      DATA_TX_PLCWI            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CARAC_PLCWI      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLCWI           : in  std_logic;                                   --! Data ready flag
      -- ppl_64_rx_sync_fsm (PLRSF) interface
      DATA_TX_PLRSF            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CARAC_PLRSF      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLRSF           : in  std_logic;                                   --! Data ready flag
      LOSS_OF_SIGNAL_PLRSF     : in  std_logic;                                   --! Loss of signal flag from PLRSF
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI      : in  std_logic;                                   --! Wait send data signal for SKIP insertion
      -- ppl_64_lane_ctrl_word_detection (PLCWD) interface
      DATA_RX_PLPL             : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CHARAC_PLPL      : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLPL            : out std_logic;                                   --! Data ready flag
      LOSS_OF_SIGNAL_PLPL      : out std_logic;                                   --! Loss of signal flag from PLPL 
      -- MIB interface
      PARALLEL_LOOPBACK_EN_MIB : in  std_logic                                    --! Enable or disable the parallel loopback
    );
  end component;

  component ppl_64_lane_init_fsm
    port (
      RST_N                               : in  std_logic;                      --! Global reset signal, Active Low
      CLK                                 : in  std_logic;                      --! Clock generated by the GTY IP
      -- Data-Link interface
      LANE_RESET_DL                       : in  std_logic;                      --! Lane reset command from the Data-Link layer
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      NO_SIGNAL_PLCWD                     : in  std_logic;                      --! Indicates that no signal is received
      RX_NEW_WORD_PLCWD                   : in  std_logic_vector(1 downto 0);   --! Indicates a new word has been received
      DETECTED_INIT1_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT1 control word has been received
      DETECTED_INIT2_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT2 control word has been received
      DETECTED_INIT3_PLCWD                : in  std_logic_vector(1 downto 0);   --! Indicates that an INIT3 control word has been received
      DETECTED_INV_INIT1_PLCWD            : in  std_logic_vector(1 downto 0);   --! Indicates that an inverted INIT1 control word has been received
      DETECTED_INV_INIT2_PLCWD            : in  std_logic_vector(1 downto 0);   --! Indicates that an inverted INIT2 control word has been received
      DETECTED_RXERR_WORD_PLCWD           : in  std_logic_vector(1 downto 0);   --! Indicates that a RXERR control word has been detected
      DETECTED_LOSS_SIGNAL_PLCWD          : in  std_logic_vector(1 downto 0);   --! Flag LOSS_SINGAL control word detected
      DETECTED_STANDBY_PLCWD              : in  std_logic_vector(1 downto 0);   --! Flag STANDBY control word detected
      COMMA_K287_RXED_PLCWD               : in  std_logic_vector(1 downto 0);   --! Flag Comma K28.7 has been received
      SEND_RXERR_PLIF                     : out std_logic_vector(1 downto 0);   --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
      INVERT_RX_BITS_PLIF                 : out std_logic;                      --! Flag to Invert rx bit received
      NO_SIGNAL_DETECTION_ENABLED_PLIF    : out std_logic;                      --! Flag to enable the no signal function
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      STANDBY_SIGNAL_X32_PLCWI            : in  std_logic;                      --! Flag STANDBY control word has been send x32
      LOST_SIGNAL_X32_PLCWI               : in  std_logic;                      --! Flag LOST_SIGNAL control word has been send x32
      SEND_INIT1_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send INIT1 control word following by 64 pseudo-random data words
      SEND_INIT2_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send control word following by 64 pseudo-random data words
      SEND_INIT3_CTRL_WORD_PLIF           : out std_logic;                      --! Flag to send control word following by 64 pseudo-random data words
      ENABLE_TRANSM_DATA_PLIF             : out std_logic;                      --! Flag to enable to send data
      SEND_32_STANDBY_CTRL_WORDS_PLIF     : out std_logic;                      --! Flag to send STANDBY control word x32
      SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF : out std_logic;                      --! Flag to send LOSS_SIGNAL control word x32
      LOST_CAUSE_PLIF                     : out std_logic_vector(01 downto 00); --! Flag to indicate the reason of the LOST_SIGNAL
      -- ppl_64_init_hssl (PLIH) interface
      RECEIVER_DISABLED_PLIF              : out std_logic;                      --! Flag to enabled RX function of HSSL IP
      CDR_PLIF                            : out std_logic;                      --! Flag to enabled CDR_PLIF function of HSSL IP
      TRANSMITTER_DISABLED_PLIF           : out std_logic;                      --! Flag to enabled TX fonction of HSSL IP
      -- PARAMETERS and STATUS (MIB interface)
      LANE_START_MIB                      : in  std_logic;                      --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART_MIB                       : in  std_logic;                      --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET_MIB                      : in  std_logic;                      --! Asserts or de-asserts LaneReset for the lane
      LANE_STATE_PLIF                     : out std_logic_vector(03 downto 00); --! Indicates the current state of the Lane Initialization state machine
      RX_ERROR_CNT_PLIF                   : out std_logic_vector(07 downto 00); --! Counter of error detected on the RX link
      RX_ERROR_OVF_PLIF                   : out std_logic                       --! Overflow flag of the RX_ERROR_CNT_PLIF
    );
  end component;

  -- RX flow
  component ppl_64_bus_split_rx
    port (
      RST_N                        : in  std_logic;                                   --! global reset
      CLK                          : in  std_logic;                                   --! Clock synchronous of the Data-link layer
      -- Data-link layer interface
      FIFO_RX_RD_EN_DL             : in  std_logic;                                   --! FIFO RX read enable flag from the Data-link layer
      DATA_RX_PLBSR                : out std_logic_vector(31 downto 0);               --! 32-bit Data parallel
      FIFO_RX_DATA_VALID_PLBSR     : out std_logic;                                   --! Flag new data
      VALID_K_CHARAC_RX_PLBSR      : out std_logic_vector(3 downto 0);                --! 4-bit valid K character
      FAR_END_CAPA_PLBSR           : out std_logic_vector(7 downto 0);                --! Capability field received in INIT3 control word
      LANE_ACTIVE_PLBSR            : out std_logic;                                   --! Lane Active flag
      -- fifo_rx_data (PLFRD) interface
      FIFO_RX_RD_EN_PLBSR          : out std_logic;                                   --! FIFO RX read enable flag
      DATA_RX_PLFRD                : in  std_logic_vector(C_DATA_WIDTH-1  downto 0);  --! 64-bit Data parallel
      FIFO_RX_DATA_VALID_PLFRD     : in  std_logic;                                   --! Flag new data
      FIFO_RX_EMPTY_PLFRD          : in  std_logic;                                   --! Flag FIFO Empty
      VALID_K_CHARAC_RX_PLFRD      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags
      DATA_RDY_RX_PLFRD            : in  std_logic_vector(1 downto 0);                --! Data valid flag
      -- ppl_64_ctrl_fifo_rx (PLCFR) interface
      FAR_END_CAPA_PLFRC           : in std_logic_vector(7 downto 0);                 --! Capability field received in INIT3 control word
      LANE_ACTIVE_PLFRC            : in std_logic                                     --! Lane Active flag
    );
  end component;

  component ppl_64_rx_wr_en_fifo
    port (
      RST_N                            : in  std_logic;                                   --! Global reset. Active Low
      CLK                              : in  std_logic;                                   --! Clock generated by HSSL IP
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      DATA_RX_PLCWD                    : in std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data from ppl_64_lane_ctrl_word_detect
      VALID_K_CHARAC_PLCWD             : in std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags from ppl_64_lane_ctrl_word_detect
      DATA_RDY_PLCWD                   : in std_logic_vector(1 downto 0);                 --! Data valid flag from ppl_64_lane_ctrl_word_detect
      -- fifo_rx_data (PLFRD) interface
      DATA_RX_PLRWEF                    : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to fifo_rx_data
      VALID_K_CHARAC_PLRWEF             : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags to fifo_rx_data
      DATA_RDY_PLRWEF                   : out std_logic_vector(1 downto 0);                --! Data valid flag to fifo_rx_data
      DATA_WR_EN_PLRWEF                 : out std_logic                                    --! Write enable flag to fifo_rx_data
    );
  end component;

  component ppl_64_lane_ctrl_word_detect
    port (
      RST_N                            : in  std_logic;                                    --! Global reset. Active Low
      CLK                              : in  std_logic;                                    --! Clock generated by HSSL IP
      -- ppl_64_lane_init_fsm (PLIF) interface
      NO_SIGNAL_PLCWD                  : out std_logic;                                    --! Flag indicating that no signal is received
      RX_NEW_WORD_PLCWD                : out std_logic_vector(1 downto 0);                 --! Flag indicating that a new word has been received
      DETECTED_INIT1_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT1 control word received
      DETECTED_INIT2_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT2 control word received
      DETECTED_INIT3_PLCWD             : out std_logic_vector(1 downto 0);                 --! Flag indicating INIT3 control word received
      DETECTED_INV_INIT1_PLCWD         : out std_logic_vector(1 downto 0);                 --! Flag indicating INV_INIT1 control word received
      DETECTED_INV_INIT2_PLCWD         : out std_logic_vector(1 downto 0);                 --! Flag indicating INV_INIT2 control word received
      DETECTED_RXERR_WORD_PLCWD        : out std_logic_vector(1 downto 0);                 --! Flag indicating RXERR control word detected
      DETECTED_LOSS_SIGNAL_PLCWD       : out std_logic_vector(1 downto 0);                 --! Flag indicating LOSS_SIGNAL control word detected
      DETECTED_STANDBY_PLCWD           : out std_logic_vector(1 downto 0);                 --! Flag indicating STANDBY control word detected
      COMMA_K287_RXED_PLCWD            : out std_logic_vector(1 downto 0);                 --! Comma K28.7 character received flag
      CAPABILITY_PLCWD                 : out std_logic_vector(15 downto 0);                --! Capability extracted from INIT3 control word: bits [31:24] and [63:56]
      SEND_RXERR_PLIF                  : in  std_logic_vector(1 downto 0);                 --! Flag to send RXERR control word to Data-Link layer when FSM exits ACTIVE_ST
      NO_SIGNAL_DETECTION_ENABLED_PLIF : in  std_logic;                                    --! Flag to enable the no-signal detection function
      ENABLE_TRANSM_DATA_PLIF          : in  std_logic;                                    --! Flag to enable the transmission of data
      -- ppl_64_parallel_loopback (PLPL) interface
      DATA_RX_PLPL                     : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data from ppl_64_parallel_loopback
      VALID_K_CHARAC_PLPL              : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags from ppl_64_parallel_loopback
      DATA_RDY_PLPL                    : in  std_logic;                                    --! Data valid flag from ppl_64_parallel_loopback
      LOSS_OF_SIGNAL_PLPL              : in  std_logic;                                    --! Loss of signal flag from ppl_64_parallel_loopback 
      -- ppl_64_rx_wr_en_fifo (PLRWEF) interface
      DATA_RX_PLCWD                    : out std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data sent to Data-Link layer
      VALID_K_CHARAC_PLCWD             : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags sent to Data-Link layer
      DATA_RDY_PLCWD                   : out std_logic_vector(1 downto 0)                  --! Data valid flag sent to Data-Link layer
    );
  end component;

  component ppl_64_rx_sync_fsm is
    port(
      RST_N                            : in  std_logic;                                    --! Global reset. Active low
      CLK                              : in  std_logic;                                    --! Clock generated by GTY IP
      -- Data-link layer interface
      LANE_RESET_DL                    : in  std_logic;                                    --! Lane reset command from Data-Link Layer.
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      DATA_RX_PLRSF                    : out std_logic_vector(C_DATA_WIDTH-1  downto 0);   --! 64-bit data to lane_ctrl_word_detect
      VALID_K_CHARAC_PLRSF             : out std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! 8-bit valid K character flags to lane_ctrl_word_detect
      DATA_RDY_PLRSF                   : out std_logic;                                    --! Data valid flag to lane_ctrl_word_detect
      LOSS_OF_SIGNAL_PLRSF             : out  std_logic;                                   --! Loss of signal flag from PLRSF
      -- ppl_64_word_alignment (PLWA) interface
      DATA_RX_PLWA                     : in  std_logic_vector(C_DATA_WIDTH-1  downto 0);   --! 64-bit data from ppl_64_word_alignment
      VALID_K_CHARAC_PLWA              : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! 8-bit valid K character flags from ppl_64_word_alignment
      INVALID_CHAR_PLWA                : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Invalid character flags from ppl_64_word_alignment
      DISPARITY_ERR_PLWA               : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Disparity error flags from ppl_64_word_alignment
      RX_WORD_IS_ALIGNED_PLWA          : in  std_logic;                                    --! RX word is aligned from ppl_64_word_alignment
      COMMA_DET_PLWA                   : in  std_logic_vector(C_K_CHAR_WIDTH-1  downto 0); --! Flag indicates that a comma is detected on the word received
      LOSS_OF_SIGNAL_PLWA              : in  std_logic;                                    --! Loss of signal flag from PLWA
      -- PARAMETERS (MIB)
      LANE_RESET                       : in  std_logic                                     --! Asserts or de-asserts LaneReset for the lane
   );
  end component;

  component ppl_64_word_alignment is
    port (
      RST_N                   : in  std_logic;                                   --! Global reset. Active low
      CLK                     : in  std_logic;                                   --! Clock generated by HSSL IP
      -- ppl_64_rx_sync_fsm (PLRSF) interface
      DATA_RX_PLWA            : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to lane_ctrl_word_detect
      VALID_K_CHARAC_PLWA     : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags to lane_ctrl_word_detect
      DATA_RDY_PLWA           : out std_logic;                                   --! Data valid flag to lane_ctrl_word_detect
      INVALID_CHAR_PLWA       : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Invalid character flags from PLWA
      DISPARITY_ERR_PLWA      : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Disparity error flags from PLWA
      RX_WORD_IS_ALIGNED_PLWA : out std_logic;                                   --! RX word is aligned from PLWA
      COMMA_DET_PLWA          : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flag indicates that a comma is detected on the word receive from PLWA
      LOSS_OF_SIGNAL_PLWA     : out  std_logic;                                   --! Loss of signal flag from PLWA
      -- HSSL IP interface
      DATA_RX_HSSL            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data from HSSL IP
      VALID_K_CHARAC_HSSL     : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags from HSSL IP
      INVALID_CHAR_HSSL       : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Invalid character flags from HSSL IP
      DISPARITY_ERR_HSSL      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Disparity error flags from HSSL IP
      RX_WORD_IS_ALIGNED_HSSL : in  std_logic;                                   --! RX word is aligned from HSSL IP
      COMMA_DET_HSSL          : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! Flag indicates that a comma is detected on the word receive
      LOSS_OF_SIGNAL_HSSL     : in  std_logic                                    --! Loss of signal flag from HSSL IP
    );
  end component;

  component FIFO_DC is
    generic (
      G_DWIDTH                : integer := 8;                                 --! Data bus FIFO length
      G_AWIDTH                : integer := 8;                                 --! Address bus FIFO length
      G_THRESHOLD_HIGH        : integer := 2**8;                              --! High threshold
      G_THRESHOLD_LOW         : integer := 0                                  --! low threshold
    );
    port (
      RST_N                   : in  std_logic;
      -- Writing port
      WR_CLK                  : in  std_logic;                                --! Clock
      WR_DATA                 : in  std_logic_vector(G_DWIDTH-1 downto 0);    --! Data write bus
      WR_DATA_EN              : in  std_logic;                                --! Write command

      -- Reading port
      RD_CLK                  : in  std_logic;                                --! Clock
      RD_DATA                 : out std_logic_vector(G_DWIDTH-1 downto 0);    --! Data read bus
      RD_DATA_EN              : in  std_logic;                                --! Read command
      RD_DATA_VLD             : out std_logic;                                --! Data valid

      -- Command port
      CMD_FLUSH               : in  std_logic;                                --! FIFO flush
      STATUS_BUSY_FLUSH       : out std_logic;                                --! FIFO is flushing

      -- Status port
      STATUS_THRESHOLD_HIGH   : out std_logic;                                --! Threshold high reached flag (sur WR_CLK)
      STATUS_THRESHOLD_LOW    : out std_logic;                                --! Threshold low reached flag (sur RD_CLK)
      STATUS_FULL             : out std_logic;                                --! Full FIFO flag (sur WR_CLK)
      STATUS_EMPTY            : out std_logic;                                --! Empty FIFO flag (sur RD_CLK)
      STATUS_LEVEL_WR         : out std_logic_vector(G_AWIDTH-1 downto 0);    --! Niveau de remplissage de la FIFO (sur WR_CLK)
      STATUS_LEVEL_RD         : out std_logic_vector(G_AWIDTH-1 downto 0)     --! Niveau de remplissage de la FIFO (sur RD_CLK)
    );
  end component;
  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- Internal signals declaration --------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------
  -- Internal signals from ppl_64_lane_init_fsm
  signal send_rxerr_plif                      : std_logic_vector(1 downto 0);
  signal invert_rx_bits_plif                  : std_logic;
  signal no_signal_detection_enabled_plif     : std_logic;
  signal send_init1_ctrl_word_plif            : std_logic;
  signal send_init2_ctrl_word_plif            : std_logic;
  signal send_init3_ctrl_word_plif            : std_logic;
  signal enable_transm_data_plif              : std_logic;
  signal send_32_standby_ctrl_words_plif      : std_logic;
  signal send_32_loss_signal_ctrl_words_plif  : std_logic;
  signal lost_cause_plif                      : std_logic_vector(01 downto 00);

  signal transmitter_disabled_plif            : std_logic;
  signal receiver_disabled_plif               : std_logic;
  signal cdr_plif                             : std_logic;

  signal lane_state_plif                      : std_logic_vector(03 downto 00);
  signal rx_error_cnt_plif                    : std_logic_vector(07 downto 00);
  signal rx_error_ovf_plif                    : std_logic;
  -------------- TX Flow --------------------------------------
  -- Internal signals from ppl_64_bus_concat_tx
  signal data_tx_plbct                        : std_logic_vector(C_DATA_WIDTH-1  downto 0);
  signal new_data_tx_plbct                    : std_logic;
  signal valid_k_charac_tx_plbct              : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal capability_tx_plbct                  : std_logic_vector(7 downto 0);
  signal lane_reset_plbct                     : std_logic;
  signal ctrl_in_plbct                        : std_logic_vector(C_DWIDTH_CTRL_TX-1 downto 0);
  signal data_plus_k_char_plbct               : std_logic_vector(71 downto 0);
  -- Internal signals from FiFo TX ctrl
  signal ctrl_in_plfic                        : std_logic_vector(C_DWIDTH_CTRL_TX-1 downto 0);
  signal data_valid_plfic                     : std_logic;
  signal capability_tx_plfic                  : std_logic_vector (7 downto 0);
  -- Internal signals from FiFo TX data
  signal data_tx_plftd                        : std_logic_vector(71 downto 00);
  signal fifo_tx_empty_plftd                  : std_logic;
  signal data_valid_plftd                     : std_logic;
   -- Internal signals from ppl_64_lane_ctrl_word_insert
  signal rd_data_en_plcwi                     : std_logic;
  signal new_data_plcwi                       : std_logic;
  signal data_tx_plcwi                        : std_logic_vector(C_DATA_WIDTH-1 downto 00);
  signal valid_k_charac_plcwi                 : std_logic_vector(C_K_CHAR_WIDTH-1 downto 00);
  signal standby_signal_x32_plcwi             : std_logic;
  signal lost_signal_x32_plcwi                : std_logic;
   -- Internal signals from skip_insertion
  signal wait_send_data_plsi                  : std_logic;
  signal data_tx_plsi                         : std_logic_vector(C_DATA_WIDTH-1 downto 00);
  signal valid_k_charac_plsi                  : std_logic_vector(C_K_CHAR_WIDTH-1 downto 00);
   -- Internal signals from parallel_loopback
  signal data_rx_plpl                         : std_logic_vector(C_DATA_WIDTH-1 downto 00);
  signal valid_k_charac_plpl                  : std_logic_vector(C_K_CHAR_WIDTH-1 downto 00);
  signal data_rdy_plpl                        : std_logic;
  signal loss_of_signal_plpl                  : std_logic;
  -------------- HSSL  ----------------------------------------
  -- HSSL instance
  signal hssl_clock_i                         : std_logic_vector(3 downto 0);
  signal clk_tx                               : std_logic;
  signal pll_pma_lock_analog_hssl             : std_logic;
  signal tx_busy_hssl                         : std_logic;
  signal rx_pma_ll_slow_locked_hssl           : std_logic;
  signal rx_pma_loss_of_signal_hssl           : std_logic;
  signal rx_busy_hssl                         : std_logic;
  signal data_rx_hssl                         : std_logic_vector(C_DATA_WIDTH-1 downto 0);
  signal valid_k_charac_hssl                  : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal invalid_char_hssl                    : std_logic_vector(C_K_CHAR_WIDTH-1  downto 0);
  signal disparity_err_hssl                   : std_logic_vector(C_K_CHAR_WIDTH-1  downto 0);
  signal rx_word_is_aligned_hssl              : std_logic;
  signal comma_det_hssl                       : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  -- inst_ppl_64_init_hssl
  signal reset_n                              : std_logic;
  signal pll_pma_pwr_up_plih                  : std_logic;
  signal tx_driver_pwrdwn_n_plih              : std_logic;
  signal pll_pma_rst_n_plih                   : std_logic;
  signal tx_rst_n_plih                        : std_logic;
  signal rx_pma_pwr_up_plih                   : std_logic;
  signal rx_pma_rst_n_plih                    : std_logic;
  signal rx_rst_n_plih                        : std_logic;
  signal hssl_reset_done_plih                 : std_logic;
  -------------- RX Flow --------------------------------------
  -- inst_ppl_64_word_alignment
  signal data_rx_plwa                         : std_logic_vector(C_DATA_WIDTH-1 downto 0);
  signal valid_k_charac_plwa                  : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal data_rdy_plwa                        : std_logic;
  signal invalid_char_plwa                    : std_logic_vector(C_K_CHAR_WIDTH-1  downto 0);
  signal disparity_err_plwa                   : std_logic_vector(C_K_CHAR_WIDTH-1  downto 0);
  signal rx_word_is_aligned_plwa              : std_logic;
  signal comma_det_plwa                       : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal loss_of_signal_plwa                  : std_logic;  
  -- Internal signals from ppl_64_rx_sync_fsm
  signal data_rx_plrsf                        : std_logic_vector(C_DATA_WIDTH-1 downto 00);
  signal valid_k_charac_plrsf                 : std_logic_vector(C_K_CHAR_WIDTH-1  downto 00);
  signal data_rdy_plrsf                       : std_logic;
  signal loss_of_signal_plrsf                 : std_logic;  
  -- Internal signals from from ppl_64_lane_ctrl_word_detect
  signal no_signal_plcwd                      : std_logic;
  signal rx_new_word_plcwd                    : std_logic_vector(1 downto 0);
  signal detected_init1_plcwd                 : std_logic_vector(1 downto 0);
  signal detected_init2_plcwd                 : std_logic_vector(1 downto 0);
  signal detected_init3_plcwd                 : std_logic_vector(1 downto 0);
  signal detected_inv_init1_plcwd             : std_logic_vector(1 downto 0);
  signal detected_inv_init2_plcwd             : std_logic_vector(1 downto 0);
  signal detected_rxerr_word_plcwd            : std_logic_vector(1 downto 0);
  signal detected_loss_signal_plcwd           : std_logic_vector(1 downto 0);
  signal detected_standby_plcwd               : std_logic_vector(1 downto 0);
  signal comma_k287_rxed_plcwd                : std_logic_vector(1 downto 0);
  signal capability_plcwd                     : std_logic_vector(15 downto 0);
  signal data_rx_plcwd                        : std_logic_vector(C_DATA_WIDTH-1 downto 0);
  signal valid_k_charac_plcwd                 : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal data_rdy_plcwd                       : std_logic_vector(1 downto 0);
  -- Internal signals from ppl_64_rx_wr_en_fifo
  signal data_rx_plrwef                        : std_logic_vector(C_DATA_WIDTH-1 downto 0);
  signal valid_k_charac_plrwef                 : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal data_rdy_plrwef                       : std_logic_vector(1 downto 0);
  signal data_wr_en_plrwef                     : std_logic;
  signal data_plus_k_char_plrwef               : std_logic_vector(73 downto 00);
  -- Internal signals from FIFO_RX data
  signal data_plus_k_char_plfrd               : std_logic_vector(73 downto 00);
  signal data_rx_plfrd                        : std_logic_vector(C_DATA_WIDTH-1 downto 0);data_rdy_rx_plfrd
  signal valid_k_charac_rx_plfrd              : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal data_rdy_rx_plfrd                    : std_logic_vector(1 downto 0);
  signal fifo_rx_data_valid_plfrd             : std_logic;
  signal fifo_rx_empty_plfrd                  : std_logic;
  -- Internal signals from FIFO_RX ctrl
  signal lane_active_capa_in_fifo_rx          : std_logic_vector(C_DWIDTH_CTRL_RX-1 downto 0);
  signal lane_active_capa_plfrc               : std_logic_vector(C_DWIDTH_CTRL_RX-1 downto 0);
  signal lane_active_plfrc                    : std_logic;
  signal far_end_capa_plfrc                   : std_logic_vector (7 downto 0);
  signal fifo_data_valid_plfrc                : std_logic;
  -- Internal signals from ppl_64_bus_split_rx
  signal fifo_rx_rd_en_plbsr                  : std_logic;
  signal far_end_capa_plbsr                   : std_logic_vector (7 downto 0);
  -- ctrl internal signals
  signal lane_reset_dl_i                      : std_logic;

begin
  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- Output assignment -------------------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------
  -- Clock and reset
  CLK_TX_OUT                 <= clk_tx;
  RST_TX_DONE                <= hssl_reset_done_plih;
  -- Data-link interface
  FIFO_RX_EMPTY              <= fifo_rx_empty_plfrd;
  FAR_END_CAPA_DL            <= far_end_capa_plbsr;
  LANE_RESET_PPL_OUT         <= lane_reset_dl_i or LANE_RESET;
  -- MIB Interface
  LANE_STATE                 <= lane_state_plif;
  RX_ERROR_CNT               <= rx_error_cnt_plif;
  RX_ERROR_OVF               <= rx_error_ovf_plif;
  LOSS_SIGNAL                <= no_signal_plcwd;
  RX_POLARITY                <= invert_rx_bits_plif;
  FAR_END_CAPA               <= far_end_capa_plbsr;

  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- Instantiation -----------------------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------

  ------------------------------------------------------------------------------
  --! Instance of ppl_64_lane_init_fsm module
  ------------------------------------------------------------------------------
  inst_lane_init_fsm : ppl_64_lane_init_fsm
    port map (
      RST_N                                => RST_TXCLK_N,
      CLK                                  => clk_tx,
      -- Data-link layer interface
      LANE_RESET_DL                        => lane_reset_dl_i,
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      NO_SIGNAL_PLCWD                      => no_signal_plcwd,
      RX_NEW_WORD_PLCWD                    => rx_new_word_plcwd,
      DETECTED_INIT1_PLCWD                 => detected_init1_plcwd,
      DETECTED_INIT2_PLCWD                 => detected_init2_plcwd,
      DETECTED_INIT3_PLCWD                 => detected_init3_plcwd,
      DETECTED_INV_INIT1_PLCWD             => detected_inv_init1_plcwd,
      DETECTED_INV_INIT2_PLCWD             => detected_inv_init2_plcwd,
      DETECTED_RXERR_WORD_PLCWD            => detected_rxerr_word_plcwd,
      DETECTED_LOSS_SIGNAL_PLCWD           => detected_loss_signal_plcwd,
      DETECTED_STANDBY_PLCWD               => detected_standby_plcwd,
      COMMA_K287_RXED_PLCWD                => comma_k287_rxed_plcwd,
      SEND_RXERR_PLIF                      => send_rxerr_plif,
      INVERT_RX_BITS_PLIF                  => invert_rx_bits_plif,
      NO_SIGNAL_DETECTION_ENABLED_PLIF     => no_signal_detection_enabled_plif,
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      STANDBY_SIGNAL_X32_PLCWI             => standby_signal_x32_plcwi,
      LOST_SIGNAL_X32_PLCWI                => lost_signal_x32_plcwi,
      SEND_INIT1_CTRL_WORD_PLIF            => send_init1_ctrl_word_plif,
      SEND_INIT2_CTRL_WORD_PLIF            => send_init2_ctrl_word_plif,
      SEND_INIT3_CTRL_WORD_PLIF            => send_init3_ctrl_word_plif,
      ENABLE_TRANSM_DATA_PLIF              => enable_transm_data_plif,
      SEND_32_STANDBY_CTRL_WORDS_PLIF      => send_32_standby_ctrl_words_plif,
      SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF  => send_32_loss_signal_ctrl_words_pliF ,
      LOST_CAUSE_PLIF                      => lost_cause_plif,
      -- ppl_64_init_hssl (PLIH) interface
      RECEIVER_DISABLED_PLIF               => receiver_disabled_plif,
      CDR_PLIF                             => cdr_plif,
      TRANSMITTER_DISABLED_PLIF            => transmitter_disabled_plif,
      -- PARAMETERS and STATUS (MIB interface)
      LANE_START_MIB                       => LANE_START,
      AUTOSTART_MIB                        => AUTOSTART,
      LANE_RESET_MIB                       => LANE_RESET,
      LANE_STATE_PLIF                      => lane_state_plif,
      RX_ERROR_CNT_PLIF                    => rx_error_cnt_plif,
      RX_ERROR_OVF_PLIF                    => rx_error_ovf_plif
    );
  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- TX Flow -----------------------------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Instance of ppl_64_bus_concat_tx module
  ------------------------------------------------------------------------------
  inst_ppl_64_bus_concat_tx: ppl_64_bus_concat_tx
    port map(
      RST_N                        => RST_N,
      CLK                          => CLK,
      -- Data-link layer interface
      DATA_TX_DL                   => DATA_TX,
      NEW_DATA_TX_DL               => NEW_DATA_TX,
      VALID_K_CHARAC_TX_DL         => VALID_K_CHARAC_TX,
      CAPABILITY_TX_DL             => CAPABILITY_TX,
      LANE_RESET_DL                => LANE_RESET,
      -- ppl_64_data_fifo_tx (PLDFT) interface
      DATA_TX_PLBCT                => data_tx_plbct,
      NEW_DATA_TX_PLBCT            => new_data_tx_plbct,
      VALID_K_CHARAC_TX_PLBCT      => valid_k_charac_tx_plbct,
      -- ppl_64_ctrl_fifo_tx (PLCFT) interface
      CAPABILITY_TX_PLBCT          => capability_tx_plbct,
      LANE_RESET_PLBCT             => lane_reset_plbct
    );
  ------------------------------------------------------------------------------
  -- Instance of TX FIFO_1MB_wrapper module
  ------------------------------------------------------------------------------
  ctrl_in_plbct       <= lane_reset_plbct & capability_tx_plbct;
  lane_reset_dl_i     <= '0'                       when lane_state_plif = "0000" else ctrl_in_plfic(8) when data_valid_plfic ='1';
  capability_tx_plfic <= ctrl_in_plfic(7 downto 0) when data_valid_plfic ='1';

  inst_fifo_in_ctrl : FIFO_DC
    generic map(
      G_DWIDTH                => C_DWIDTH_CTRL_TX,
      G_AWIDTH                => C_AWIDTH_CTRL_TX,
      G_THRESHOLD_HIGH        => 2**C_AWIDTH_CTRL_TX,
      G_THRESHOLD_LOW         => 0
   )
    port map(
      RST_N                   => RST_TXCLK_N,
      -- Writing port
      WR_CLK                  => CLK,
      WR_DATA                 => ctrl_in_plbct,
      WR_DATA_EN              => '1',
      -- Reading port
      RD_CLK                  => clk_tx,
      RD_DATA                 => ctrl_in_plfic,
      RD_DATA_EN              => '1',
      RD_DATA_VLD             => data_valid_plfic,
      -- Command port
      CMD_FLUSH               => '0',
      STATUS_BUSY_FLUSH       => open,
      -- Status port
      STATUS_THRESHOLD_HIGH   => open,
      STATUS_THRESHOLD_LOW    => open,
      STATUS_FULL             => open,
      STATUS_EMPTY            => open,
      STATUS_LEVEL_WR         => open,
      STATUS_LEVEL_RD         => open
   );
  ------------------------------------------------------------------------------
  -- Instance of TX FIFO_1MB_wrapper module
  ------------------------------------------------------------------------------
  data_plus_k_char_plbct   <= valid_k_charac_tx_plbct & data_tx_plbct;

  inst_fifo_tx_data : FIFO_DC
  generic map(
       G_DWIDTH                => C_DWIDTH,
       G_AWIDTH                => C_AWIDTH_TX,
       G_THRESHOLD_HIGH        => 2**C_AWIDTH_TX,
       G_THRESHOLD_LOW         => 0
   )
   port map(
       RST_N                   => RST_TXCLK_N,
       -- Writing port
       WR_CLK                  => CLK,
       WR_DATA                 => data_plus_k_char_plbct,
       WR_DATA_EN              => new_data_tx_plbct,
       -- Reading port
       RD_CLK                  => clk_tx,
       RD_DATA                 => data_tx_plftd,
       RD_DATA_EN              => rd_data_en_plcwi,
       RD_DATA_VLD             => data_valid_plftd,
       -- Command port
       CMD_FLUSH               => LANE_RESET_DL,
       STATUS_BUSY_FLUSH       => open,
       -- Status port
       STATUS_THRESHOLD_HIGH   => open,
       STATUS_THRESHOLD_LOW    => open,
       STATUS_FULL             => FIFO_TX_FULL,
       STATUS_EMPTY            => fifo_tx_empty_plftd,
       STATUS_LEVEL_WR         => open,
       STATUS_LEVEL_RD         => open
   );

  ------------------------------------------------------------------------------
  -- Instance of ppl_64_lane_ctrl_word_insert module
  ------------------------------------------------------------------------------
  inst_ppl_64_lane_ctrl_word_insert: ppl_64_lane_ctrl_word_insert
    port map(
      RST_N                                => RST_TXCLK_N,
      CLK                                  => clk_tx,
      -- Data-Link interface
      RD_DATA_EN_PLCWI                     => rd_data_en_plcwi,
      RD_DATA_VALID_DL                     => data_valid_plftd,
      CAPABILITY_DL                        => capability_tx_plfic,
      DATA_TX_DL                           => data_tx_plftd(63 downto 0),
      VALID_K_CHARAC_DL                    => data_tx_plftd(71 downto 64),
      NO_DATA_DL                           => fifo_tx_empty_plftd,
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI                  => wait_send_data_plsi,
      NEW_DATA_PLCWI                       => new_data_plcwi,
      DATA_TX_PLCWI                        => data_tx_plcwi,
      VALID_K_CHARAC_PLCWI                 => valid_k_charac_plcwi,
      -- ppl_64_lane_init_fsm (PLIF) interface
      SEND_INIT1_CTRL_WORD_PLIF            => send_init1_ctrl_word_plif,
      SEND_INIT2_CTRL_WORD_PLIF            => send_init2_ctrl_word_plif,
      SEND_INIT3_CTRL_WORD_PLIF            => send_init3_ctrl_word_plif,
      ENABLE_TRANSM_DATA_PLIF              => enable_transm_data_plif,
      SEND_32_STANDBY_CTRL_WORDS_PLIF      => send_32_standby_ctrl_words_plif,
      SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF  => send_32_loss_signal_ctrl_words_plif,
      STANDBY_SIGNAL_X32_PLCWI             => standby_signal_x32_plcwi,
      LOST_SIGNAL_X32_PLCWI                => lost_signal_x32_plcwi,
      LOST_CAUSE_PLIF                      => lost_cause_plif,
      -- MIB interface
      STANDBY_REASON_MIB                   => STANDBY_REASON

   );

  ------------------------------------------------------------------------------
  -- Instance of skip_insertion module
  ------------------------------------------------------------------------------
  inst_ppl_64_skip_insertion: ppl_64_skip_insertion
    port map (
      RST_N                   => RST_TXCLK_N,
      CLK                     => clk_tx,
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      NEW_DATA_PLCWI          => new_data_plcwi,
      DATA_TX_PLCWI           => data_tx_plcwi,
      VALID_K_CHARAC_PLCWI    => valid_k_charac_plcwi,
      WAIT_SEND_DATA_PLSI     => wait_send_data_plsi,
      -- HSSL interface
      DATA_TX_PLSI            => data_tx_plsi,
      VALID_K_CHARAC_PLSI     => valid_k_charac_plsi,
      -- ppl_64_lane_init_fsm (PLIF) interface
      ENABLE_TRANSM_DATA_PLIF => enable_transm_data_plif
    );

  ------------------------------------------------------------------------------
  -- Instance of parallel_loopback module
  ------------------------------------------------------------------------------
  inst_ppl_64_parallel_loopback : ppl_64_parallel_loopback
    port map(
      CLK                      => RST_TXCLK_N,
      RST_N                    => clk_tx,
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      DATA_TX_PLCWI            => data_tx_plcwi,
      VALID_K_CARAC_PLCWI      => valid_k_charac_plcwi,
      DATA_RDY_PLCWI           => new_data_plcwi,
      -- ppl_64_rx_sync_fsm (PLRSF) interface
      DATA_TX_PLRSF            => data_rx_plrsf,
      VALID_K_CARAC_PLRSF      => valid_k_charac_plrsf,
      DATA_RDY_PLRSF           => data_rdy_plrsf,
      LOSS_OF_SIGNAL_PLRSF     => loss_of_signal_plrsf,
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI      => wait_send_data_plsi,
      --ppl_64_lane_ctrl_word_detection (PLCWD) interface
      DATA_RX_PLPL             => data_rx_plpl,
      VALID_K_CHARAC_PLPL      => valid_k_charac_plpl,
      DATA_RDY_PLPL            => data_rdy_plpl,
      LOSS_OF_SIGNAL_PLPL      => loss_of_signal_plpl,
      -- MIB interface
      PARALLEL_LOOPBACK_EN_MIB => parallel_loopback_en
    );
  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- HSSL --------------------------------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------
  hssl_clock_i(0) <= clk_tx;
  hssl_clock_i(1) <= clk_tx;
  hssl_clock_i(2) <= clk_tx;
  hssl_clock_i(3) <= clk_tx;
  ------------------------------------------------------------------------------
  -- Instance of hssl module
  ------------------------------------------------------------------------------
  inst_SpaceFibre_64b : SpaceFibre_64b
    port map (
      HSSL_CLOCK_I                => hssl_clock_i,
      RX0N                        => RX_NEG,
      RX0P                        => RX_POS,
      RX1N                        => '1',
      RX1P                        => '0',
      RX2N                        => '1',
      RX2P                        => '0',
      RX3N                        => '1',
      RX3P                        => '0',
      TX0N                        => TX_NEG,
      TX0P                        => TX_POS,
      TX1N                        => open,
      TX1P                        => open,
      TX2N                        => open,
      TX2P                        => open,
      TX3N                        => open,
      TX3P                        => open,
      CKREFN                      => CLK_REF_N,
      CKREFP                      => CLK_REF_P,
      CLOCK_O                     => clk_tx,
      DYN_CFG_EN_I                => '0',
      DYN_ADDR_I                  => (others => '0'),
      DYN_CALIBRATION_CS_N_I      => '1',
      DYN_LANE_CS_N_I             => "1111",
      DYN_WDATA_I                 => (others => '0'),
      DYN_WDATA_SEL_I             => '0',
      DYN_WE_N_I                  => '1',
      PLL_PMA_LOCK_ANALOG         => pll_pma_lock_analog_hssl,
      PLL_PMA_PWR_UP_I            => pll_pma_pwr_up_plih,
      PLL_PMA_RST_N_I             => pll_pma_rst_n_plih,
      PLL_LOCK                    => open,
      TX0_BUSY_O                  => tx_busy_hssl,
      TX0_CLK_ENA_I               => '1',
      TX0_CLK_O                   => open,
      TX0_DATA_I                  => data_tx_plsi,
      TX0_CTRL_DRIVER_PWRDWN_N_I  => tx_driver_pwrdwn_n_plih,
      TX0_RST_N_I                 => tx_rst_n_plih,
      TX0_CTRL_CHAR_IS_K_I        => valid_k_charac_plsi,
      RX0_BUSY_O                  => rx_busy_hssl,
      RX0_CTRL_EL_BUFF_STAT_O     => open,
      RX0_CTRL_CHAR_IS_ALIGNED_O  => rx_word_is_aligned_hssl,
      RX0_CTRL_CHAR_IS_COMMA_O    => comma_det_hssl,
      RX0_CTRL_CHAR_IS_F_O        => open,
      RX0_CTRL_CHAR_IS_K_O        => valid_k_charac_hssl,
      RX0_CTRL_DISP_ERR_O         => disparity_err_hssl,
      RX0_CTRL_NOT_IN_TABLE_O     => invalid_char_hssl,
      RX0_CTRL_VALID_REALIGN_O    => open,
      RX0_DATA_O                  => data_rx_hssl,
      RX0_OVS_BIT_SEL_I           => "00",
      RX0_EYE_RST_I               => '0',
      RX0_PMA_LL_FAST_LOCKED_O    => open,
      RX0_PMA_LL_SLOW_LOCKED_O    => rx_pma_ll_slow_locked_hssl,
      RX0_PMA_LOSS_OF_SIGNAL_O    => rx_pma_loss_of_signal_hssl,
      RX0_PMA_PLL_LOCK_O          => open,
      RX0_PMA_PLL_LOCK_TRACK_O    => open,
      RX0_PMA_RST_N_I             => rx_pma_rst_n_plih,
      RX0_PMA_PWR_UP_I            => rx_pma_pwr_up_plih,
      RX0_RST_N_I                 => rx_rst_n_plih,
      RX0_TEST_O                  => open,
      RX0_REPLACE_EN_I            => '0',
      RX0_ALIGN_SYNC_I            => '1',
      RX0_EL_BUFF_RST_I           => '0'
    );
  ------------------------------------------------------------------------------
  -- Instance of ppl_64_init_hssl module
  ------------------------------------------------------------------------------
  reset_n <= RST_N and not(LANE_RESET) and not(lane_reset_dl_i);

  inst_ppl_64_init_hssl: ppl_64_init_hssl
    port map (
      RST_N                      => reset_n,
      CLK                        => CLK,
      -- ppl_64_lane_init_fsm (PLIF) interface
      RECEIVER_DISABLED_PLIF     => receiver_disabled_plif,
      CDR_PLIF                   => cdr_plif,
      TRANSMITTER_DISABLED_PLIF  => transmitter_disabled_plif,
      -- HSSL interface
      PLL_PMA_PWR_UP_PLIH        => pll_pma_pwr_up_plih,
      TX_DRIVER_PWRDWN_N_PLIH    => tx_driver_pwrdwn_n_plih,
      PLL_PMA_RST_N_PLIH         => pll_pma_rst_n_plih,
      PLL_PMA_LOCK_ANALOG_HSSL   => pll_pma_lock_analog_hssl,
      TX_RST_N_PLIH              => tx_rst_n_plih,
      TX_BUSY_HSSL               => tx_busy_hssl,
      RX_PMA_PWR_UP_PLIH         => rx_pma_pwr_up_plih,
      RX_PMA_RST_N_PLIH          => rx_pma_rst_n_plih,
      RX_PMA_LL_SLOW_LOCKED_HSSL => rx_pma_ll_slow_locked_hssl,
      RX_RST_N_PLIH              => rx_rst_n_plih,
      RX_BUSY_HSSL               => rx_busy_hssl,
      -- Output
      HSSL_RESET_DONE_PLIH       => hssl_reset_done_plih
  );
  ----------------------------------------------------------------------------------------------------------------------------------------
  -------------------------------------------------------- RX Flow -----------------------------------------------------------------------
  ----------------------------------------------------------------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Instance of ppl_64_word_alignment module
  ------------------------------------------------------------------------------
  inst_ppl_64_word_alignment : ppl_64_word_alignment
    port map(
      RST_N                   => RST_TXCLK_N,
      CLK                     => clk_tx,
      -- ppl_64_rx_sync_fsm (PLRSF) interface
      DATA_RX_PLWA            => data_rx_plwa,
      VALID_K_CHARAC_PLWA     => valid_k_charac_plwa,
      DATA_RDY_PLWA           => data_rdy_plwa,
      INVALID_CHAR_PLWA       => invalid_char_plwa,
      DISPARITY_ERR_PLWA      => disparity_err_plwa,
      RX_WORD_IS_ALIGNED_PLWA => rx_word_is_aligned_plwa,
      COMMA_DET_PLWA          => comma_det_plwa,
      LOSS_OF_SIGNAL_PLWA     => loss_of_signal_plwa,
      -- HSSL IP interface
      DATA_RX_HSSL            => data_rx_hssl,
      VALID_K_CHARAC_HSSL     => valid_k_charac_hssl,
      INVALID_CHAR_HSSL       => invalid_char_hssl,
      DISPARITY_ERR_HSSL      => disparity_err_hssl,
      RX_WORD_IS_ALIGNED_HSSL => rx_word_is_aligned_hssl,
      COMMA_DET_HSSL          => comma_det_hssl,
      LOSS_OF_SIGNAL_HSSL     => rx_pma_loss_of_signal_hssl
    );
  ------------------------------------------------------------------------------
  -- Instance of rx_sync_fsm module
  ------------------------------------------------------------------------------
  inst_ppl_64_rx_sync_fsm : ppl_64_rx_sync_fsm
    port map(
      RST_N                   => RST_TXCLK_N,
      CLK                     => clk_tx,
      -- Data-link layer interface
      LANE_RESET_DL           => LANE_RESET_DL,
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      DATA_RX_PLRSF           => data_rx_plrsf,
      VALID_K_CHARAC_PLRSF    => valid_k_charac_plrsf,
      DATA_RDY_PLRSF          => data_rdy_plrsf,
      LOSS_OF_SIGNAL_PLRSF    => loss_of_signal_plrsf,
      -- ppl_64_word_alignment (PLWA) interface
      DATA_RX_PLWA            => data_rx_plwa,
      VALID_K_CHARAC_PLWA     => valid_k_charac_plwa,
      INVALID_CHAR_PLWA       => invalid_char_plwa,
      DISPARITY_ERR_PLWA      => disparity_err_plwa,
      RX_WORD_IS_ALIGNED_PLWA => rx_word_is_aligned_plwa,
      COMMA_DET_PLWA          => comma_det_plwa,
      LOSS_OF_SIGNAL_PLWA     => loss_of_signal_plwa,
      -- PARAMETERS (MIB)
      LANE_RESET              => lane_reset
    );

  ------------------------------------------------------------------------------
  -- Instance of ppl_64_lane_ctrl_word_detect module
  ------------------------------------------------------------------------------
  inst_lane_ctrl_word_detect : ppl_64_lane_ctrl_word_detect
    port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- ppl_64_lane_init_fsm (PLIF) interface
      NO_SIGNAL_PLCWD                  => no_signal_plcwd,
      RX_NEW_WORD_PLCWD                => rx_new_word_plcwd,
      DETECTED_INIT1_PLCWD             => detected_init1_plcwd,
      DETECTED_INIT2_PLCWD             => detected_init2_plcwd,
      DETECTED_INIT3_PLCWD             => detected_init3_plcwd,
      DETECTED_INV_INIT1_PLCWD         => detected_inv_init1_plcwd,
      DETECTED_INV_INIT2_PLCWD         => detected_inv_init2_plcwd,
      DETECTED_RXERR_WORD_PLCWD        => detected_rxerr_word_plcwd,
      DETECTED_LOSS_SIGNAL_PLCWD       => detected_loss_signal_plcwd,
      DETECTED_STANDBY_PLCWD           => detected_standby_plcwd,
      COMMA_K287_RXED_PLCWD            => comma_k287_rxed_plcwd,
      CAPABILITY_PLCWD                 => capability_plcwd,
      SEND_RXERR_PLIF                  => send_rxerr_plif,
      NO_SIGNAL_DETECTION_ENABLED_PLIF => no_signal_detection_enabled_plif,
      ENABLE_TRANSM_DATA_PLIF          => enable_transm_data_plif,
      -- ppl_64_parallel_loopback (PLPL) interface
      DATA_RX_PLPL                     => data_rx_plpl,
      VALID_K_CHARAC_PLPL              => valid_k_charac_plpl,
      DATA_RDY_PLPL                    => data_rdy_plpl,
      LOSS_OF_SIGNAL_PLPL              => loss_of_signal_plpl,
      -- ppl_64_rx_wr_en_fifo (PLRWEF) interface
      DATA_RX_PLCWD                    => data_rx_plcwd,
      VALID_K_CHARAC_PLCWD             => valid_k_charac_plcwd,
      DATA_RDY_PLCWD                   => data_rdy_plcwd
  );

  ------------------------------------------------------------------------------
  -- Instance of ppl_64_rx_wr_en_fifo module
  ------------------------------------------------------------------------------
  inst_ppl_64_rx_wr_en_fifo: ppl_64_rx_wr_en_fifo
    port map(
      RST_N                            => RST_TXCLK_N,
      CLK                              => clk_tx,
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      DATA_RX_PLCWD                    => data_rx_plcwd,
      VALID_K_CHARAC_PLCWD             => valid_k_charac_plcwd,
      DATA_RDY_PLCWD                   => data_rdy_plcwd,
      -- fifo_rx_data (PLFRD) interface
      DATA_RX_PLRWEF                    => data_rx_plrwef,
      VALID_K_CHARAC_PLRWEF             => valid_k_charac_plrwef,
      DATA_RDY_PLRWEF                   => data_rdy_plrwef,
      DATA_WR_EN_PLRWEF                 => data_wr_en_plrwef
    );
  ------------------------------------------------------------------------------
  -- Instance of RX FIFO_1MB_wrapper module
  ------------------------------------------------------------------------------
  data_plus_k_char_plrwef   <= data_rdy_plrwef & valid_k_charac_plrwef & data_rx_plrwef;   -- regroup data and valid K char and ready on 74-bit vector

  inst_fifo_rx_data : FIFO_DC
     generic map(
          G_DWIDTH                => C_DWIDTH + C_RDY_WORD,
          G_AWIDTH                => C_AWIDTH_RX,
          G_THRESHOLD_HIGH        => 2**C_AWIDTH_RX,
          G_THRESHOLD_LOW         => 0
      )
      port map(
          RST_N                   => RST_N,
          -- Writing port
          WR_CLK                  => clk_tx,
          WR_DATA                 => data_plus_k_char_plrwef,
          WR_DATA_EN              => data_wr_en_plrwef,
          -- Reading port
          RD_CLK                  => CLK,
          RD_DATA                 => data_plus_k_char_plfrd,
          RD_DATA_EN              => fifo_rx_rd_en_plbsr,
          RD_DATA_VLD             => fifo_rx_data_valid_plfrd,
          -- Command port
          CMD_FLUSH               => LANE_RESET_DL,
          STATUS_BUSY_FLUSH       => open,
          -- Status port
          STATUS_THRESHOLD_HIGH   => open,
          STATUS_THRESHOLD_LOW    => open,
          STATUS_FULL             => open,
          STATUS_EMPTY            => fifo_rx_empty_plfrd,
          STATUS_LEVEL_WR         => open,
          STATUS_LEVEL_RD         => open
      );
  ------------------------------------------------------------------------------
  -- Instance of TX FIFO_1MB_wrapper module
  ------------------------------------------------------------------------------
  lane_active_capa_in_fifo_rx <= enable_transm_data_plif & capability_plcwd(15 downto 8);
  lane_active_plfrc           <= lane_active_capa_plfrc(8)          when fifo_data_valid_plfrc ='1';
  far_end_capa_plfrc          <= lane_active_capa_plfrc(7 downto 0) when fifo_data_valid_plfrc ='1';
  inst_fifo_rx_ctrl : FIFO_DC
  generic map(
       G_DWIDTH                => C_DWIDTH_CTRL_RX,
       G_AWIDTH                => C_AWIDTH_CTRL_RX,
       G_THRESHOLD_HIGH        => 2**C_AWIDTH_CTRL_RX,
       G_THRESHOLD_LOW         => 0
   )
   port map(
       RST_N                   => RST_N,
       -- Writing port
       WR_CLK                  => clk_tx,
       WR_DATA                 => lane_active_capa_in_fifo_rx,
       WR_DATA_EN              => '1',
       -- Reading port
       RD_CLK                  => CLK,
       RD_DATA                 => lane_active_capa_plfrc,
       RD_DATA_EN              => '1',
       RD_DATA_VLD             => fifo_data_valid_plfrc,
       -- Command port
       CMD_FLUSH               => '0',
       STATUS_BUSY_FLUSH       => open,
       -- Status port
       STATUS_THRESHOLD_HIGH   => open,
       STATUS_THRESHOLD_LOW    => open,
       STATUS_FULL             => open,
       STATUS_EMPTY            => open,
       STATUS_LEVEL_WR         => open,
       STATUS_LEVEL_RD         => open
   );
  ------------------------------------------------------------------------------
  -- Instance of ppl_64_bus_split_rx
  ------------------------------------------------------------------------------
  data_rx_plfrd           <= data_plus_k_char_plfrd (63 downto 0);
  valid_k_charac_rx_plfrd <= data_plus_k_char_plfrd (71 downto 64);
  data_rdy_rx_plfrd       <= data_plus_k_char_plfrd (73 downto 72);
  inst_ppl_64_bus_split_rx : ppl_64_bus_split_rx
    port map (
      RST_N                       => RST_N,
      CLK                         => CLK,
      -- Data-link layer interface
      FIFO_RX_RD_EN_DL            => FIFO_RX_RD_EN,
      DATA_RX_PLBSR               => DATA_RX,
      FIFO_RX_DATA_VALID_PLBSR    => FIFO_RX_DATA_VALID,
      VALID_K_CHARAC_RX_PLBSR     => VALID_K_CHARAC_RX,
      FAR_END_CAPA_PLBSR          => far_end_capa_plbsr,
      LANE_ACTIVE_PLBSR           => LANE_ACTIVE_DL,
      -- fifo_rx_data (PLFRD) interface
      FIFO_RX_RD_EN_PLBSR         => fifo_rx_rd_en_plbsr,
      DATA_RX_PLFRD               => data_rx_plfrd,
      FIFO_RX_DATA_VALID_PLFRD    => fifo_rx_data_valid_plfrd,
      FIFO_RX_EMPTY_PLFRD         => fifo_rx_empty_plfrd,
      VALID_K_CHARAC_RX_PLFRD     => valid_k_charac_rx_plfrd,
      DATA_RDY_RX_PLFRD           => data_rdy_rx_plfrd,
      -- ppl_64_ctrl_fifo_rx (PLCFR) interface
      FAR_END_CAPA_PLFRC          => far_end_capa_plfrc,
      LANE_ACTIVE_PLFRC           => lane_active_plfrc
    );

end architecture rtl;
