// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_VCU_DEFINES_VH
`else
`define B_VCU_DEFINES_VH

// Look-up table parameters
//

`define VCU_ADDR_N  15
`define VCU_ADDR_SZ 32
`define VCU_DATA_SZ 40

// Attribute addresses
//

`define VCU__CORECLKREQ    32'h0000
`define VCU__CORECLKREQ_SZ 32

`define VCU__DECHORRESOLUTION    32'h0001
`define VCU__DECHORRESOLUTION_SZ 32

`define VCU__DECODERCHROMAFORMAT    32'h0002
`define VCU__DECODERCHROMAFORMAT_SZ 40

`define VCU__DECODERCODING    32'h0003
`define VCU__DECODERCODING_SZ 40

`define VCU__DECODERCOLORDEPTH    32'h0004
`define VCU__DECODERCOLORDEPTH_SZ 32

`define VCU__DECODERNUMCORES    32'h0005
`define VCU__DECODERNUMCORES_SZ 32

`define VCU__DECVERTRESOLUTION    32'h0006
`define VCU__DECVERTRESOLUTION_SZ 32

`define VCU__ENABLEDECODER    32'h0007
`define VCU__ENABLEDECODER_SZ 40

`define VCU__ENABLEENCODER    32'h0008
`define VCU__ENABLEENCODER_SZ 40

`define VCU__ENCHORRESOLUTION    32'h0009
`define VCU__ENCHORRESOLUTION_SZ 32

`define VCU__ENCODERCHROMAFORMAT    32'h000a
`define VCU__ENCODERCHROMAFORMAT_SZ 40

`define VCU__ENCODERCODING    32'h000b
`define VCU__ENCODERCODING_SZ 40

`define VCU__ENCODERCOLORDEPTH    32'h000c
`define VCU__ENCODERCOLORDEPTH_SZ 32

`define VCU__ENCODERNUMCORES    32'h000d
`define VCU__ENCODERNUMCORES_SZ 32

`define VCU__ENCVERTRESOLUTION    32'h000e
`define VCU__ENCVERTRESOLUTION_SZ 32

`endif  // B_VCU_DEFINES_VH