// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_MBUFGCE_DIV_DEFINES_VH
`else
`define B_MBUFGCE_DIV_DEFINES_VH

// Look-up table parameters
//

`define MBUFGCE_DIV_ADDR_N  8
`define MBUFGCE_DIV_ADDR_SZ 32
`define MBUFGCE_DIV_DATA_SZ 88

// Attribute addresses
//

`define MBUFGCE_DIV__BUFGCE_DIVIDE    32'h00000000
`define MBUFGCE_DIV__BUFGCE_DIVIDE_SZ 32

`define MBUFGCE_DIV__CE_TYPE    32'h00000001
`define MBUFGCE_DIV__CE_TYPE_SZ 64

`define MBUFGCE_DIV__HARDSYNC_CLR    32'h00000002
`define MBUFGCE_DIV__HARDSYNC_CLR_SZ 40

`define MBUFGCE_DIV__IS_CE_INVERTED    32'h00000003
`define MBUFGCE_DIV__IS_CE_INVERTED_SZ 1

`define MBUFGCE_DIV__IS_CLR_INVERTED    32'h00000004
`define MBUFGCE_DIV__IS_CLR_INVERTED_SZ 1

`define MBUFGCE_DIV__IS_I_INVERTED    32'h00000005
`define MBUFGCE_DIV__IS_I_INVERTED_SZ 1

`define MBUFGCE_DIV__MODE    32'h00000006
`define MBUFGCE_DIV__MODE_SZ 88

`define MBUFGCE_DIV__STARTUP_SYNC    32'h00000007
`define MBUFGCE_DIV__STARTUP_SYNC_SZ 40

`endif  // B_MBUFGCE_DIV_DEFINES_VH