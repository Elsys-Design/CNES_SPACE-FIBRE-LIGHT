// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_PCIE40E5_DEFINES_VH
`else
`define B_PCIE40E5_DEFINES_VH

// Look-up table parameters
//

`define PCIE40E5_ADDR_N  756
`define PCIE40E5_ADDR_SZ 32
`define PCIE40E5_DATA_SZ 144

// Attribute addresses
//

`define PCIE40E5__AER_CAP_PERMIT_ROOTERR_UPDATE    32'h00000000
`define PCIE40E5__AER_CAP_PERMIT_ROOTERR_UPDATE_SZ 40

`define PCIE40E5__ARI_CAP_ENABLE    32'h00000001
`define PCIE40E5__ARI_CAP_ENABLE_SZ 40

`define PCIE40E5__AUTO_FLR_RESPONSE    32'h00000002
`define PCIE40E5__AUTO_FLR_RESPONSE_SZ 40

`define PCIE40E5__AXISTEN_IF_CCIX_RX_CREDIT_LIMIT    32'h00000003
`define PCIE40E5__AXISTEN_IF_CCIX_RX_CREDIT_LIMIT_SZ 8

`define PCIE40E5__AXISTEN_IF_CCIX_TX_CREDIT_LIMIT    32'h00000004
`define PCIE40E5__AXISTEN_IF_CCIX_TX_CREDIT_LIMIT_SZ 6

`define PCIE40E5__AXISTEN_IF_CCIX_TX_REGISTERED_TREADY    32'h00000005
`define PCIE40E5__AXISTEN_IF_CCIX_TX_REGISTERED_TREADY_SZ 40

`define PCIE40E5__AXISTEN_IF_CC_ALIGNMENT_MODE    32'h00000006
`define PCIE40E5__AXISTEN_IF_CC_ALIGNMENT_MODE_SZ 2

`define PCIE40E5__AXISTEN_IF_COMPL_TIMEOUT_REG0    32'h00000007
`define PCIE40E5__AXISTEN_IF_COMPL_TIMEOUT_REG0_SZ 24

`define PCIE40E5__AXISTEN_IF_COMPL_TIMEOUT_REG1    32'h00000008
`define PCIE40E5__AXISTEN_IF_COMPL_TIMEOUT_REG1_SZ 28

`define PCIE40E5__AXISTEN_IF_CQ_ALIGNMENT_MODE    32'h00000009
`define PCIE40E5__AXISTEN_IF_CQ_ALIGNMENT_MODE_SZ 2

`define PCIE40E5__AXISTEN_IF_CQ_EN_POISONED_MEM_WR    32'h0000000a
`define PCIE40E5__AXISTEN_IF_CQ_EN_POISONED_MEM_WR_SZ 40

`define PCIE40E5__AXISTEN_IF_CQ_POISON_DISCARD_DISABLE    32'h0000000b
`define PCIE40E5__AXISTEN_IF_CQ_POISON_DISCARD_DISABLE_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_10B_TAGS    32'h0000000c
`define PCIE40E5__AXISTEN_IF_ENABLE_10B_TAGS_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_256_TAGS    32'h0000000d
`define PCIE40E5__AXISTEN_IF_ENABLE_256_TAGS_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_CLIENT_TAG    32'h0000000e
`define PCIE40E5__AXISTEN_IF_ENABLE_CLIENT_TAG_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE    32'h0000000f
`define PCIE40E5__AXISTEN_IF_ENABLE_INTERNAL_MSIX_TABLE_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK    32'h00000010
`define PCIE40E5__AXISTEN_IF_ENABLE_MESSAGE_RID_CHECK_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_MSG_ROUTE    32'h00000011
`define PCIE40E5__AXISTEN_IF_ENABLE_MSG_ROUTE_SZ 18

`define PCIE40E5__AXISTEN_IF_ENABLE_RX_MSG_INTFC    32'h00000012
`define PCIE40E5__AXISTEN_IF_ENABLE_RX_MSG_INTFC_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_RX_TAG_SCALING    32'h00000013
`define PCIE40E5__AXISTEN_IF_ENABLE_RX_TAG_SCALING_SZ 40

`define PCIE40E5__AXISTEN_IF_ENABLE_TX_TAG_SCALING    32'h00000014
`define PCIE40E5__AXISTEN_IF_ENABLE_TX_TAG_SCALING_SZ 40

`define PCIE40E5__AXISTEN_IF_EXTEND_CPL_TIMEOUT    32'h00000015
`define PCIE40E5__AXISTEN_IF_EXTEND_CPL_TIMEOUT_SZ 2

`define PCIE40E5__AXISTEN_IF_EXT_512    32'h00000016
`define PCIE40E5__AXISTEN_IF_EXT_512_SZ 40

`define PCIE40E5__AXISTEN_IF_EXT_512_CC_STRADDLE    32'h00000017
`define PCIE40E5__AXISTEN_IF_EXT_512_CC_STRADDLE_SZ 40

`define PCIE40E5__AXISTEN_IF_EXT_512_CQ_STRADDLE    32'h00000018
`define PCIE40E5__AXISTEN_IF_EXT_512_CQ_STRADDLE_SZ 40

`define PCIE40E5__AXISTEN_IF_EXT_512_RC_STRADDLE    32'h00000019
`define PCIE40E5__AXISTEN_IF_EXT_512_RC_STRADDLE_SZ 40

`define PCIE40E5__AXISTEN_IF_EXT_512_RQ_STRADDLE    32'h0000001a
`define PCIE40E5__AXISTEN_IF_EXT_512_RQ_STRADDLE_SZ 40

`define PCIE40E5__AXISTEN_IF_INTERNAL_MSIX_VECTORS_PER_FUNCTION    32'h0000001b
`define PCIE40E5__AXISTEN_IF_INTERNAL_MSIX_VECTORS_PER_FUNCTION_SZ 2

`define PCIE40E5__AXISTEN_IF_LEGACY_MODE_ENABLE    32'h0000001c
`define PCIE40E5__AXISTEN_IF_LEGACY_MODE_ENABLE_SZ 40

`define PCIE40E5__AXISTEN_IF_MSIX_FROM_RAM_PIPELINE    32'h0000001d
`define PCIE40E5__AXISTEN_IF_MSIX_FROM_RAM_PIPELINE_SZ 40

`define PCIE40E5__AXISTEN_IF_MSIX_RX_PARITY_EN    32'h0000001e
`define PCIE40E5__AXISTEN_IF_MSIX_RX_PARITY_EN_SZ 40

`define PCIE40E5__AXISTEN_IF_MSIX_TO_RAM_PIPELINE    32'h0000001f
`define PCIE40E5__AXISTEN_IF_MSIX_TO_RAM_PIPELINE_SZ 40

`define PCIE40E5__AXISTEN_IF_PASID_UR_CHECK_DISABLE    32'h00000020
`define PCIE40E5__AXISTEN_IF_PASID_UR_CHECK_DISABLE_SZ 40

`define PCIE40E5__AXISTEN_IF_RC_ALIGNMENT_MODE    32'h00000021
`define PCIE40E5__AXISTEN_IF_RC_ALIGNMENT_MODE_SZ 2

`define PCIE40E5__AXISTEN_IF_RC_STRADDLE    32'h00000022
`define PCIE40E5__AXISTEN_IF_RC_STRADDLE_SZ 40

`define PCIE40E5__AXISTEN_IF_RQ_ALIGNMENT_MODE    32'h00000023
`define PCIE40E5__AXISTEN_IF_RQ_ALIGNMENT_MODE_SZ 2

`define PCIE40E5__AXISTEN_IF_RQ_CC_REGISTERED_TREADY    32'h00000024
`define PCIE40E5__AXISTEN_IF_RQ_CC_REGISTERED_TREADY_SZ 40

`define PCIE40E5__AXISTEN_IF_RX_PARITY_EN    32'h00000025
`define PCIE40E5__AXISTEN_IF_RX_PARITY_EN_SZ 40

`define PCIE40E5__AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT    32'h00000026
`define PCIE40E5__AXISTEN_IF_SIM_SHORT_CPL_TIMEOUT_SZ 40

`define PCIE40E5__AXISTEN_IF_TX_PARITY_EN    32'h00000027
`define PCIE40E5__AXISTEN_IF_TX_PARITY_EN_SZ 40

`define PCIE40E5__AXISTEN_IF_WIDTH    32'h00000028
`define PCIE40E5__AXISTEN_IF_WIDTH_SZ 2

`define PCIE40E5__AXISTEN_USER_SPARE    32'h00000029
`define PCIE40E5__AXISTEN_USER_SPARE_SZ 16

`define PCIE40E5__CCIX_CFG_MGMT_MUX_ENABLE    32'h0000002a
`define PCIE40E5__CCIX_CFG_MGMT_MUX_ENABLE_SZ 40

`define PCIE40E5__CCIX_DIRECT_ATTACH_MODE    32'h0000002b
`define PCIE40E5__CCIX_DIRECT_ATTACH_MODE_SZ 40

`define PCIE40E5__CCIX_ENABLE    32'h0000002c
`define PCIE40E5__CCIX_ENABLE_SZ 40

`define PCIE40E5__CCIX_OPT_TLP_GEN_AND_RECEPT_EN_CONTROL_INTERNAL    32'h0000002d
`define PCIE40E5__CCIX_OPT_TLP_GEN_AND_RECEPT_EN_CONTROL_INTERNAL_SZ 40

`define PCIE40E5__CCIX_PDVSEC_CPL_TIMEOUT    32'h0000002e
`define PCIE40E5__CCIX_PDVSEC_CPL_TIMEOUT_SZ 17

`define PCIE40E5__CCIX_PROTOCOL_PF0_DVSEC_ENABLE    32'h0000002f
`define PCIE40E5__CCIX_PROTOCOL_PF0_DVSEC_ENABLE_SZ 40

`define PCIE40E5__CCIX_PROTOCOL_PF1_DVSEC_ENABLE    32'h00000030
`define PCIE40E5__CCIX_PROTOCOL_PF1_DVSEC_ENABLE_SZ 40

`define PCIE40E5__CCIX_TRANSPORT_PF0_DVSEC_ENABLE    32'h00000031
`define PCIE40E5__CCIX_TRANSPORT_PF0_DVSEC_ENABLE_SZ 40

`define PCIE40E5__CCIX_TX_CREDIT_CHECK_DISABLE    32'h00000032
`define PCIE40E5__CCIX_TX_CREDIT_CHECK_DISABLE_SZ 40

`define PCIE40E5__CCIX_VENDOR_ID    32'h00000033
`define PCIE40E5__CCIX_VENDOR_ID_SZ 16

`define PCIE40E5__CFG_BYPASS_MODE_ENABLE    32'h00000034
`define PCIE40E5__CFG_BYPASS_MODE_ENABLE_SZ 40

`define PCIE40E5__CFG_PRIVATE_SPC    32'h00000035
`define PCIE40E5__CFG_PRIVATE_SPC_SZ 40

`define PCIE40E5__CFG_SPEC_4_0    32'h00000036
`define PCIE40E5__CFG_SPEC_4_0_SZ 40

`define PCIE40E5__CRM_CORE_CLK_FREQ    32'h00000037
`define PCIE40E5__CRM_CORE_CLK_FREQ_SZ 5

`define PCIE40E5__CRM_USER_CLK_FREQ    32'h00000038
`define PCIE40E5__CRM_USER_CLK_FREQ_SZ 3

`define PCIE40E5__DEBUG_AXI4ST_SPARE    32'h00000039
`define PCIE40E5__DEBUG_AXI4ST_SPARE_SZ 16

`define PCIE40E5__DEBUG_AXIST_DISABLE_FEATURE_BIT    32'h0000003a
`define PCIE40E5__DEBUG_AXIST_DISABLE_FEATURE_BIT_SZ 8

`define PCIE40E5__DEBUG_CAR_SPARE    32'h0000003b
`define PCIE40E5__DEBUG_CAR_SPARE_SZ 4

`define PCIE40E5__DEBUG_CFG_SPARE    32'h0000003c
`define PCIE40E5__DEBUG_CFG_SPARE_SZ 16

`define PCIE40E5__DEBUG_LL_SPARE    32'h0000003d
`define PCIE40E5__DEBUG_LL_SPARE_SZ 16

`define PCIE40E5__DEBUG_NO_STICKY_RESET    32'h0000003e
`define PCIE40E5__DEBUG_NO_STICKY_RESET_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR    32'h0000003f
`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_DEFRAMER_ERROR_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR    32'h00000040
`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_ERROR_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR    32'h00000041
`define PCIE40E5__DEBUG_PL_DISABLE_LES_UPDATE_ON_SKP_PARITY_ERROR_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL    32'h00000042
`define PCIE40E5__DEBUG_PL_DISABLE_REC_ENTRY_ON_DYNAMIC_DSKEW_FAIL_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW    32'h00000043
`define PCIE40E5__DEBUG_PL_DISABLE_REC_ENTRY_ON_RX_BUFFER_UNDER_OVER_FLOW_SZ 40

`define PCIE40E5__DEBUG_PL_DISABLE_SCRAMBLING    32'h00000044
`define PCIE40E5__DEBUG_PL_DISABLE_SCRAMBLING_SZ 40

`define PCIE40E5__DEBUG_PL_SIM_RESET_LFSR    32'h00000045
`define PCIE40E5__DEBUG_PL_SIM_RESET_LFSR_SZ 40

`define PCIE40E5__DEBUG_PL_SPARE    32'h00000046
`define PCIE40E5__DEBUG_PL_SPARE_SZ 16

`define PCIE40E5__DEBUG_TL_DISABLE_FC_TIMEOUT    32'h00000047
`define PCIE40E5__DEBUG_TL_DISABLE_FC_TIMEOUT_SZ 40

`define PCIE40E5__DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS    32'h00000048
`define PCIE40E5__DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_SZ 40

`define PCIE40E5__DEBUG_TL_SPARE    32'h00000049
`define PCIE40E5__DEBUG_TL_SPARE_SZ 16

`define PCIE40E5__DELAYED_FLR    32'h0000004a
`define PCIE40E5__DELAYED_FLR_SZ 40

`define PCIE40E5__DNSTREAM_LINK_NUM    32'h0000004b
`define PCIE40E5__DNSTREAM_LINK_NUM_SZ 8

`define PCIE40E5__DSN_CAP_ENABLE    32'h0000004c
`define PCIE40E5__DSN_CAP_ENABLE_SZ 40

`define PCIE40E5__EXTENDED_CFG_EXTEND_INTERFACE_ENABLE    32'h0000004d
`define PCIE40E5__EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_SZ 40

`define PCIE40E5__HEADER_TYPE_OVERRIDE    32'h0000004e
`define PCIE40E5__HEADER_TYPE_OVERRIDE_SZ 40

`define PCIE40E5__IS_SWITCH_PORT    32'h0000004f
`define PCIE40E5__IS_SWITCH_PORT_SZ 40

`define PCIE40E5__LEGACY_CFG_EXTEND_INTERFACE_ENABLE    32'h00000050
`define PCIE40E5__LEGACY_CFG_EXTEND_INTERFACE_ENABLE_SZ 40

`define PCIE40E5__LINK_CONTROL2_SELECTABLE_DEEMPH    32'h00000051
`define PCIE40E5__LINK_CONTROL2_SELECTABLE_DEEMPH_SZ 40

`define PCIE40E5__LL_ACK_TIMEOUT    32'h00000052
`define PCIE40E5__LL_ACK_TIMEOUT_SZ 9

`define PCIE40E5__LL_ACK_TIMEOUT_EN    32'h00000053
`define PCIE40E5__LL_ACK_TIMEOUT_EN_SZ 40

`define PCIE40E5__LL_ACK_TIMEOUT_FUNC    32'h00000054
`define PCIE40E5__LL_ACK_TIMEOUT_FUNC_SZ 2

`define PCIE40E5__LL_DISABLE_SCHED_TX_NAK    32'h00000055
`define PCIE40E5__LL_DISABLE_SCHED_TX_NAK_SZ 40

`define PCIE40E5__LL_FEATURE_EN_DLLP_EXCHANGE    32'h00000056
`define PCIE40E5__LL_FEATURE_EN_DLLP_EXCHANGE_SZ 40

`define PCIE40E5__LL_FEATURE_EN_FC_SCALING    32'h00000057
`define PCIE40E5__LL_FEATURE_EN_FC_SCALING_SZ 40

`define PCIE40E5__LL_FEATURE_EN_FC_SCALING_SCALE_FACTOR_4    32'h00000058
`define PCIE40E5__LL_FEATURE_EN_FC_SCALING_SCALE_FACTOR_4_SZ 40

`define PCIE40E5__LL_REPLAY_FROM_RAM_PIPELINE    32'h00000059
`define PCIE40E5__LL_REPLAY_FROM_RAM_PIPELINE_SZ 40

`define PCIE40E5__LL_REPLAY_TIMEOUT    32'h0000005a
`define PCIE40E5__LL_REPLAY_TIMEOUT_SZ 9

`define PCIE40E5__LL_REPLAY_TIMEOUT_EN    32'h0000005b
`define PCIE40E5__LL_REPLAY_TIMEOUT_EN_SZ 40

`define PCIE40E5__LL_REPLAY_TIMEOUT_FUNC    32'h0000005c
`define PCIE40E5__LL_REPLAY_TIMEOUT_FUNC_SZ 2

`define PCIE40E5__LL_REPLAY_TIMER40_ENABLE    32'h0000005d
`define PCIE40E5__LL_REPLAY_TIMER40_ENABLE_SZ 40

`define PCIE40E5__LL_REPLAY_TO_RAM_PIPELINE    32'h0000005e
`define PCIE40E5__LL_REPLAY_TO_RAM_PIPELINE_SZ 40

`define PCIE40E5__LL_RX_TLP_PARITY_GEN    32'h0000005f
`define PCIE40E5__LL_RX_TLP_PARITY_GEN_SZ 40

`define PCIE40E5__LL_TX_PARITY_CHECK_CHANGE_DISABLE    32'h00000060
`define PCIE40E5__LL_TX_PARITY_CHECK_CHANGE_DISABLE_SZ 40

`define PCIE40E5__LL_TX_STALL_ON_ASPM_L1_ENTRY_DISABLE    32'h00000061
`define PCIE40E5__LL_TX_STALL_ON_ASPM_L1_ENTRY_DISABLE_SZ 40

`define PCIE40E5__LL_TX_STALL_ON_PPM_L1_ENTRY_DISABLE    32'h00000062
`define PCIE40E5__LL_TX_STALL_ON_PPM_L1_ENTRY_DISABLE_SZ 40

`define PCIE40E5__LL_TX_TLP_PARITY_CHK    32'h00000063
`define PCIE40E5__LL_TX_TLP_PARITY_CHK_SZ 40

`define PCIE40E5__LL_UFC_ARBITER_ENABLE    32'h00000064
`define PCIE40E5__LL_UFC_ARBITER_ENABLE_SZ 40

`define PCIE40E5__LL_USER_SPARE    32'h00000065
`define PCIE40E5__LL_USER_SPARE_SZ 16

`define PCIE40E5__LTR_TX_MESSAGE_MINIMUM_INTERVAL    32'h00000066
`define PCIE40E5__LTR_TX_MESSAGE_MINIMUM_INTERVAL_SZ 10

`define PCIE40E5__LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE    32'h00000067
`define PCIE40E5__LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_SZ 40

`define PCIE40E5__LTR_TX_MESSAGE_ON_LTR_ENABLE    32'h00000068
`define PCIE40E5__LTR_TX_MESSAGE_ON_LTR_ENABLE_SZ 40

`define PCIE40E5__MCAP_CAP_NEXTPTR    32'h00000069
`define PCIE40E5__MCAP_CAP_NEXTPTR_SZ 12

`define PCIE40E5__MCAP_CFG_SLAVE_BLOCK    32'h0000006a
`define PCIE40E5__MCAP_CFG_SLAVE_BLOCK_SZ 40

`define PCIE40E5__MCAP_CONFIGURE_OVERRIDE    32'h0000006b
`define PCIE40E5__MCAP_CONFIGURE_OVERRIDE_SZ 40

`define PCIE40E5__MCAP_ENABLE    32'h0000006c
`define PCIE40E5__MCAP_ENABLE_SZ 40

`define PCIE40E5__MCAP_EOS_DESIGN_SWITCH    32'h0000006d
`define PCIE40E5__MCAP_EOS_DESIGN_SWITCH_SZ 40

`define PCIE40E5__MCAP_FPGA_BITSTREAM_VERSION    32'h0000006e
`define PCIE40E5__MCAP_FPGA_BITSTREAM_VERSION_SZ 32

`define PCIE40E5__MCAP_GATE_IO_ENABLE_DESIGN_SWITCH    32'h0000006f
`define PCIE40E5__MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_SZ 40

`define PCIE40E5__MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH    32'h00000070
`define PCIE40E5__MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_SZ 40

`define PCIE40E5__MCAP_INPUT_GATE_DESIGN_SWITCH    32'h00000071
`define PCIE40E5__MCAP_INPUT_GATE_DESIGN_SWITCH_SZ 40

`define PCIE40E5__MCAP_INTERRUPT_ON_MCAP_EOS    32'h00000072
`define PCIE40E5__MCAP_INTERRUPT_ON_MCAP_EOS_SZ 40

`define PCIE40E5__MCAP_INTERRUPT_ON_MCAP_ERROR    32'h00000073
`define PCIE40E5__MCAP_INTERRUPT_ON_MCAP_ERROR_SZ 40

`define PCIE40E5__MCAP_VSEC_ID    32'h00000074
`define PCIE40E5__MCAP_VSEC_ID_SZ 16

`define PCIE40E5__MCAP_VSEC_LEN    32'h00000075
`define PCIE40E5__MCAP_VSEC_LEN_SZ 12

`define PCIE40E5__MCAP_VSEC_REV    32'h00000076
`define PCIE40E5__MCAP_VSEC_REV_SZ 4

`define PCIE40E5__PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE    32'h00000077
`define PCIE40E5__PF0_AER_CAP_ECRC_GEN_AND_CHECK_CAPABLE_SZ 40

`define PCIE40E5__PF0_AER_CAP_NEXTPTR    32'h00000078
`define PCIE40E5__PF0_AER_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_ARI_CAP_NEXTPTR    32'h00000079
`define PCIE40E5__PF0_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_ARI_CAP_NEXT_FUNC    32'h0000007a
`define PCIE40E5__PF0_ARI_CAP_NEXT_FUNC_SZ 8

`define PCIE40E5__PF0_ARI_CAP_VER    32'h0000007b
`define PCIE40E5__PF0_ARI_CAP_VER_SZ 4

`define PCIE40E5__PF0_ATS_CAP_INV_QUEUE_DEPTH    32'h0000007c
`define PCIE40E5__PF0_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__PF0_ATS_CAP_NEXTPTR    32'h0000007d
`define PCIE40E5__PF0_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_ATS_CAP_ON    32'h0000007e
`define PCIE40E5__PF0_ATS_CAP_ON_SZ 40

`define PCIE40E5__PF0_BAR0_APERTURE_SIZE    32'h0000007f
`define PCIE40E5__PF0_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_BAR0_CONTROL    32'h00000080
`define PCIE40E5__PF0_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF0_BAR1_APERTURE_SIZE    32'h00000081
`define PCIE40E5__PF0_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_BAR1_CONTROL    32'h00000082
`define PCIE40E5__PF0_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF0_BAR2_APERTURE_SIZE    32'h00000083
`define PCIE40E5__PF0_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_BAR2_CONTROL    32'h00000084
`define PCIE40E5__PF0_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF0_BAR3_APERTURE_SIZE    32'h00000085
`define PCIE40E5__PF0_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_BAR3_CONTROL    32'h00000086
`define PCIE40E5__PF0_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF0_BAR4_APERTURE_SIZE    32'h00000087
`define PCIE40E5__PF0_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_BAR4_CONTROL    32'h00000088
`define PCIE40E5__PF0_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF0_BAR5_APERTURE_SIZE    32'h00000089
`define PCIE40E5__PF0_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_BAR5_CONTROL    32'h0000008a
`define PCIE40E5__PF0_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF0_CAPABILITY_POINTER    32'h0000008b
`define PCIE40E5__PF0_CAPABILITY_POINTER_SZ 8

`define PCIE40E5__PF0_CCIX_ESM_QUICK_EQ_TIMEOUT    32'h0000008c
`define PCIE40E5__PF0_CCIX_ESM_QUICK_EQ_TIMEOUT_SZ 3

`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_ID    32'h0000008d
`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_ID_SZ 16

`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_LENGTH    32'h0000008e
`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_LENGTH_SZ 12

`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_NEXTPTR    32'h0000008f
`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_REVISION    32'h00000090
`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_REVISION_SZ 4

`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_VENDOR_ID    32'h00000091
`define PCIE40E5__PF0_CCIX_PDVSEC_CAP_VENDOR_ID_SZ 16

`define PCIE40E5__PF0_CCIX_PDVSEC_PCR_SIZE    32'h00000092
`define PCIE40E5__PF0_CCIX_PDVSEC_PCR_SIZE_SZ 12

`define PCIE40E5__PF0_CCIX_PDVSEC_PCR_START_ADDR    32'h00000093
`define PCIE40E5__PF0_CCIX_PDVSEC_PCR_START_ADDR_SZ 12

`define PCIE40E5__PF0_CCIX_PDVSEC_PCSR_SIZE    32'h00000094
`define PCIE40E5__PF0_CCIX_PDVSEC_PCSR_SIZE_SZ 12

`define PCIE40E5__PF0_CCIX_PDVSEC_PCSR_START_ADDR    32'h00000095
`define PCIE40E5__PF0_CCIX_PDVSEC_PCSR_START_ADDR_SZ 12

`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_ID    32'h00000096
`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_ID_SZ 16

`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_LENGTH    32'h00000097
`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_LENGTH_SZ 12

`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_NEXTPTR    32'h00000098
`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_REVISION    32'h00000099
`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_REVISION_SZ 4

`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_VENDOR_ID    32'h0000009a
`define PCIE40E5__PF0_CCIX_TDVSEC_CAP_VENDOR_ID_SZ 16

`define PCIE40E5__PF0_CCIX_TDVSEC_CCIX_VC_BYTE_OFFSET    32'h0000009b
`define PCIE40E5__PF0_CCIX_TDVSEC_CCIX_VC_BYTE_OFFSET_SZ 7

`define PCIE40E5__PF0_CLASS_CODE    32'h0000009c
`define PCIE40E5__PF0_CLASS_CODE_SZ 24

`define PCIE40E5__PF0_DEV_CAP2_10B_TAG_COMPLETER_SUPPORTED    32'h0000009d
`define PCIE40E5__PF0_DEV_CAP2_10B_TAG_COMPLETER_SUPPORTED_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_10B_TAG_REQUESTER_SUPPORTED    32'h0000009e
`define PCIE40E5__PF0_DEV_CAP2_10B_TAG_REQUESTER_SUPPORTED_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT    32'h0000009f
`define PCIE40E5__PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT    32'h000000a0
`define PCIE40E5__PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT    32'h000000a1
`define PCIE40E5__PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_ARI_FORWARD_ENABLE    32'h000000a2
`define PCIE40E5__PF0_DEV_CAP2_ARI_FORWARD_ENABLE_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE    32'h000000a3
`define PCIE40E5__PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_LTR_SUPPORT    32'h000000a4
`define PCIE40E5__PF0_DEV_CAP2_LTR_SUPPORT_SZ 40

`define PCIE40E5__PF0_DEV_CAP2_OBFF_SUPPORT    32'h000000a5
`define PCIE40E5__PF0_DEV_CAP2_OBFF_SUPPORT_SZ 2

`define PCIE40E5__PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT    32'h000000a6
`define PCIE40E5__PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_SZ 40

`define PCIE40E5__PF0_DEV_CAP_ENDPOINT_L0S_LATENCY    32'h000000a7
`define PCIE40E5__PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_SZ 3

`define PCIE40E5__PF0_DEV_CAP_ENDPOINT_L1_LATENCY    32'h000000a8
`define PCIE40E5__PF0_DEV_CAP_ENDPOINT_L1_LATENCY_SZ 3

`define PCIE40E5__PF0_DEV_CAP_EXT_TAG_SUPPORTED    32'h000000a9
`define PCIE40E5__PF0_DEV_CAP_EXT_TAG_SUPPORTED_SZ 40

`define PCIE40E5__PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE    32'h000000aa
`define PCIE40E5__PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_SZ 40

`define PCIE40E5__PF0_DEV_CAP_MAX_PAYLOAD_SIZE    32'h000000ab
`define PCIE40E5__PF0_DEV_CAP_MAX_PAYLOAD_SIZE_SZ 3

`define PCIE40E5__PF0_DEV_CONTROL2_PERMIT_IDO_CPL_EN    32'h000000ac
`define PCIE40E5__PF0_DEV_CONTROL2_PERMIT_IDO_CPL_EN_SZ 40

`define PCIE40E5__PF0_DEV_CONTROL2_PERMIT_IDO_REQ_EN    32'h000000ad
`define PCIE40E5__PF0_DEV_CONTROL2_PERMIT_IDO_REQ_EN_SZ 40

`define PCIE40E5__PF0_DLL_FEATURE_CAP_ID    32'h000000ae
`define PCIE40E5__PF0_DLL_FEATURE_CAP_ID_SZ 16

`define PCIE40E5__PF0_DLL_FEATURE_CAP_NEXTPTR    32'h000000af
`define PCIE40E5__PF0_DLL_FEATURE_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_DLL_FEATURE_CAP_ON    32'h000000b0
`define PCIE40E5__PF0_DLL_FEATURE_CAP_ON_SZ 40

`define PCIE40E5__PF0_DLL_FEATURE_CAP_VER    32'h000000b1
`define PCIE40E5__PF0_DLL_FEATURE_CAP_VER_SZ 4

`define PCIE40E5__PF0_DSN_CAP_NEXTPTR    32'h000000b2
`define PCIE40E5__PF0_DSN_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_EXPANSION_ROM_APERTURE_SIZE    32'h000000b3
`define PCIE40E5__PF0_EXPANSION_ROM_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_EXPANSION_ROM_ENABLE    32'h000000b4
`define PCIE40E5__PF0_EXPANSION_ROM_ENABLE_SZ 40

`define PCIE40E5__PF0_INTERRUPT_PIN    32'h000000b5
`define PCIE40E5__PF0_INTERRUPT_PIN_SZ 3

`define PCIE40E5__PF0_LINK_CAP_ASPM_SUPPORT    32'h000000b6
`define PCIE40E5__PF0_LINK_CAP_ASPM_SUPPORT_SZ 2

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    32'h000000b7
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    32'h000000b8
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3    32'h000000b9
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4    32'h000000ba
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN4_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1    32'h000000bb
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2    32'h000000bc
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3    32'h000000bd
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4    32'h000000be
`define PCIE40E5__PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN4_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1    32'h000000bf
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2    32'h000000c0
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3    32'h000000c1
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4    32'h000000c2
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN4_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1    32'h000000c3
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2    32'h000000c4
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3    32'h000000c5
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_SZ 3

`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4    32'h000000c6
`define PCIE40E5__PF0_LINK_CAP_L1_EXIT_LATENCY_GEN4_SZ 3

`define PCIE40E5__PF0_LINK_CONTROL_RCB    32'h000000c7
`define PCIE40E5__PF0_LINK_CONTROL_RCB_SZ 1

`define PCIE40E5__PF0_LINK_STATUS_SLOT_CLOCK_CONFIG    32'h000000c8
`define PCIE40E5__PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_SZ 40

`define PCIE40E5__PF0_LTR_CAP_MAX_NOSNOOP_LAT    32'h000000c9
`define PCIE40E5__PF0_LTR_CAP_MAX_NOSNOOP_LAT_SZ 10

`define PCIE40E5__PF0_LTR_CAP_MAX_SNOOP_LAT    32'h000000ca
`define PCIE40E5__PF0_LTR_CAP_MAX_SNOOP_LAT_SZ 10

`define PCIE40E5__PF0_LTR_CAP_NEXTPTR    32'h000000cb
`define PCIE40E5__PF0_LTR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_LTR_CAP_VER    32'h000000cc
`define PCIE40E5__PF0_LTR_CAP_VER_SZ 4

`define PCIE40E5__PF0_MARGINING_CAP_ID    32'h000000cd
`define PCIE40E5__PF0_MARGINING_CAP_ID_SZ 16

`define PCIE40E5__PF0_MARGINING_CAP_NEXTPTR    32'h000000ce
`define PCIE40E5__PF0_MARGINING_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_MARGINING_CAP_ON    32'h000000cf
`define PCIE40E5__PF0_MARGINING_CAP_ON_SZ 40

`define PCIE40E5__PF0_MARGINING_CAP_VER    32'h000000d0
`define PCIE40E5__PF0_MARGINING_CAP_VER_SZ 4

`define PCIE40E5__PF0_MARGINING_USES_DRVR_SW    32'h000000d1
`define PCIE40E5__PF0_MARGINING_USES_DRVR_SW_SZ 40

`define PCIE40E5__PF0_MSIX_CAP_NEXTPTR    32'h000000d2
`define PCIE40E5__PF0_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF0_MSIX_CAP_PBA_BIR    32'h000000d3
`define PCIE40E5__PF0_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__PF0_MSIX_CAP_PBA_OFFSET    32'h000000d4
`define PCIE40E5__PF0_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__PF0_MSIX_CAP_TABLE_BIR    32'h000000d5
`define PCIE40E5__PF0_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__PF0_MSIX_CAP_TABLE_OFFSET    32'h000000d6
`define PCIE40E5__PF0_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__PF0_MSIX_CAP_TABLE_SIZE    32'h000000d7
`define PCIE40E5__PF0_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__PF0_MSIX_VECTOR_COUNT    32'h000000d8
`define PCIE40E5__PF0_MSIX_VECTOR_COUNT_SZ 6

`define PCIE40E5__PF0_MSI_CAP_MULTIMSGCAP    32'h000000d9
`define PCIE40E5__PF0_MSI_CAP_MULTIMSGCAP_SZ 3

`define PCIE40E5__PF0_MSI_CAP_NEXTPTR    32'h000000da
`define PCIE40E5__PF0_MSI_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF0_MSI_CAP_PERVECMASKCAP    32'h000000db
`define PCIE40E5__PF0_MSI_CAP_PERVECMASKCAP_SZ 40

`define PCIE40E5__PF0_PASID_CAP_EXEC_PERM_SUPP    32'h000000dc
`define PCIE40E5__PF0_PASID_CAP_EXEC_PERM_SUPP_SZ 1

`define PCIE40E5__PF0_PASID_CAP_MAX_PASID_WIDTH    32'h000000dd
`define PCIE40E5__PF0_PASID_CAP_MAX_PASID_WIDTH_SZ 5

`define PCIE40E5__PF0_PASID_CAP_NEXTPTR    32'h000000de
`define PCIE40E5__PF0_PASID_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_PASID_CAP_ON    32'h000000df
`define PCIE40E5__PF0_PASID_CAP_ON_SZ 1

`define PCIE40E5__PF0_PASID_CAP_PRIVIL_MODE_SUPP    32'h000000e0
`define PCIE40E5__PF0_PASID_CAP_PRIVIL_MODE_SUPP_SZ 1

`define PCIE40E5__PF0_PCIE_CAP_NEXTPTR    32'h000000e1
`define PCIE40E5__PF0_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF0_PL16_CAP_ID    32'h000000e2
`define PCIE40E5__PF0_PL16_CAP_ID_SZ 16

`define PCIE40E5__PF0_PL16_CAP_NEXTPTR    32'h000000e3
`define PCIE40E5__PF0_PL16_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_PL16_CAP_ON    32'h000000e4
`define PCIE40E5__PF0_PL16_CAP_ON_SZ 40

`define PCIE40E5__PF0_PL16_CAP_VER    32'h000000e5
`define PCIE40E5__PF0_PL16_CAP_VER_SZ 4

`define PCIE40E5__PF0_PM_CAP_ID    32'h000000e6
`define PCIE40E5__PF0_PM_CAP_ID_SZ 8

`define PCIE40E5__PF0_PM_CAP_NEXTPTR    32'h000000e7
`define PCIE40E5__PF0_PM_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D0    32'h000000e8
`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D0_SZ 40

`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D1    32'h000000e9
`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D1_SZ 40

`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D3COLD    32'h000000ea
`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D3COLD_SZ 40

`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D3HOT    32'h000000eb
`define PCIE40E5__PF0_PM_CAP_PMESUPPORT_D3HOT_SZ 40

`define PCIE40E5__PF0_PM_CAP_SUPP_D1_STATE    32'h000000ec
`define PCIE40E5__PF0_PM_CAP_SUPP_D1_STATE_SZ 40

`define PCIE40E5__PF0_PM_CAP_VER_ID    32'h000000ed
`define PCIE40E5__PF0_PM_CAP_VER_ID_SZ 3

`define PCIE40E5__PF0_PM_CSR_NOSOFTRESET    32'h000000ee
`define PCIE40E5__PF0_PM_CSR_NOSOFTRESET_SZ 40

`define PCIE40E5__PF0_PRI_CAP_NEXTPTR    32'h000000ef
`define PCIE40E5__PF0_PRI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_PRI_CAP_ON    32'h000000f0
`define PCIE40E5__PF0_PRI_CAP_ON_SZ 40

`define PCIE40E5__PF0_PRI_OST_PR_CAPACITY    32'h000000f1
`define PCIE40E5__PF0_PRI_OST_PR_CAPACITY_SZ 32

`define PCIE40E5__PF0_SECONDARY_PCIE_CAP_NEXTPTR    32'h000000f2
`define PCIE40E5__PF0_SECONDARY_PCIE_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED    32'h000000f3
`define PCIE40E5__PF0_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ 40

`define PCIE40E5__PF0_SRIOV_BAR0_APERTURE_SIZE    32'h000000f4
`define PCIE40E5__PF0_SRIOV_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_SRIOV_BAR0_CONTROL    32'h000000f5
`define PCIE40E5__PF0_SRIOV_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_BAR1_APERTURE_SIZE    32'h000000f6
`define PCIE40E5__PF0_SRIOV_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_SRIOV_BAR1_CONTROL    32'h000000f7
`define PCIE40E5__PF0_SRIOV_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_BAR2_APERTURE_SIZE    32'h000000f8
`define PCIE40E5__PF0_SRIOV_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_SRIOV_BAR2_CONTROL    32'h000000f9
`define PCIE40E5__PF0_SRIOV_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_BAR3_APERTURE_SIZE    32'h000000fa
`define PCIE40E5__PF0_SRIOV_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_SRIOV_BAR3_CONTROL    32'h000000fb
`define PCIE40E5__PF0_SRIOV_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_BAR4_APERTURE_SIZE    32'h000000fc
`define PCIE40E5__PF0_SRIOV_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF0_SRIOV_BAR4_CONTROL    32'h000000fd
`define PCIE40E5__PF0_SRIOV_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_BAR5_APERTURE_SIZE    32'h000000fe
`define PCIE40E5__PF0_SRIOV_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF0_SRIOV_BAR5_CONTROL    32'h000000ff
`define PCIE40E5__PF0_SRIOV_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF0_SRIOV_CAP_INITIAL_VF    32'h00000100
`define PCIE40E5__PF0_SRIOV_CAP_INITIAL_VF_SZ 16

`define PCIE40E5__PF0_SRIOV_CAP_NEXTPTR    32'h00000101
`define PCIE40E5__PF0_SRIOV_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_SRIOV_CAP_TOTAL_VF    32'h00000102
`define PCIE40E5__PF0_SRIOV_CAP_TOTAL_VF_SZ 16

`define PCIE40E5__PF0_SRIOV_CAP_VER    32'h00000103
`define PCIE40E5__PF0_SRIOV_CAP_VER_SZ 4

`define PCIE40E5__PF0_SRIOV_FIRST_VF_OFFSET    32'h00000104
`define PCIE40E5__PF0_SRIOV_FIRST_VF_OFFSET_SZ 16

`define PCIE40E5__PF0_SRIOV_FUNC_DEP_LINK    32'h00000105
`define PCIE40E5__PF0_SRIOV_FUNC_DEP_LINK_SZ 16

`define PCIE40E5__PF0_SRIOV_SUPPORTED_PAGE_SIZE    32'h00000106
`define PCIE40E5__PF0_SRIOV_SUPPORTED_PAGE_SIZE_SZ 32

`define PCIE40E5__PF0_SRIOV_VF_DEVICE_ID    32'h00000107
`define PCIE40E5__PF0_SRIOV_VF_DEVICE_ID_SZ 16

`define PCIE40E5__PF0_TPHR_CAP_DEV_SPECIFIC_MODE    32'h00000108
`define PCIE40E5__PF0_TPHR_CAP_DEV_SPECIFIC_MODE_SZ 40

`define PCIE40E5__PF0_TPHR_CAP_ENABLE    32'h00000109
`define PCIE40E5__PF0_TPHR_CAP_ENABLE_SZ 40

`define PCIE40E5__PF0_TPHR_CAP_INT_VEC_MODE    32'h0000010a
`define PCIE40E5__PF0_TPHR_CAP_INT_VEC_MODE_SZ 40

`define PCIE40E5__PF0_TPHR_CAP_NEXTPTR    32'h0000010b
`define PCIE40E5__PF0_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_TPHR_CAP_ST_MODE_SEL    32'h0000010c
`define PCIE40E5__PF0_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__PF0_TPHR_CAP_ST_TABLE_LOC    32'h0000010d
`define PCIE40E5__PF0_TPHR_CAP_ST_TABLE_LOC_SZ 2

`define PCIE40E5__PF0_TPHR_CAP_ST_TABLE_SIZE    32'h0000010e
`define PCIE40E5__PF0_TPHR_CAP_ST_TABLE_SIZE_SZ 11

`define PCIE40E5__PF0_TPHR_CAP_VER    32'h0000010f
`define PCIE40E5__PF0_TPHR_CAP_VER_SZ 4

`define PCIE40E5__PF0_VC_ARB_CAPABILITY    32'h00000110
`define PCIE40E5__PF0_VC_ARB_CAPABILITY_SZ 4

`define PCIE40E5__PF0_VC_ARB_TBL_OFFSET    32'h00000111
`define PCIE40E5__PF0_VC_ARB_TBL_OFFSET_SZ 8

`define PCIE40E5__PF0_VC_CAP_ENABLE    32'h00000112
`define PCIE40E5__PF0_VC_CAP_ENABLE_SZ 40

`define PCIE40E5__PF0_VC_CAP_NEXTPTR    32'h00000113
`define PCIE40E5__PF0_VC_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF0_VC_CAP_VER    32'h00000114
`define PCIE40E5__PF0_VC_CAP_VER_SZ 4

`define PCIE40E5__PF0_VC_EXTENDED_COUNT    32'h00000115
`define PCIE40E5__PF0_VC_EXTENDED_COUNT_SZ 40

`define PCIE40E5__PF0_VC_LOW_PRIORITY_EXTENDED_COUNT    32'h00000116
`define PCIE40E5__PF0_VC_LOW_PRIORITY_EXTENDED_COUNT_SZ 40

`define PCIE40E5__PF1_AER_CAP_NEXTPTR    32'h00000117
`define PCIE40E5__PF1_AER_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_ARI_CAP_NEXTPTR    32'h00000118
`define PCIE40E5__PF1_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_ARI_CAP_NEXT_FUNC    32'h00000119
`define PCIE40E5__PF1_ARI_CAP_NEXT_FUNC_SZ 8

`define PCIE40E5__PF1_ATS_CAP_INV_QUEUE_DEPTH    32'h0000011a
`define PCIE40E5__PF1_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__PF1_ATS_CAP_NEXTPTR    32'h0000011b
`define PCIE40E5__PF1_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_ATS_CAP_ON    32'h0000011c
`define PCIE40E5__PF1_ATS_CAP_ON_SZ 40

`define PCIE40E5__PF1_BAR0_APERTURE_SIZE    32'h0000011d
`define PCIE40E5__PF1_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_BAR0_CONTROL    32'h0000011e
`define PCIE40E5__PF1_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF1_BAR1_APERTURE_SIZE    32'h0000011f
`define PCIE40E5__PF1_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_BAR1_CONTROL    32'h00000120
`define PCIE40E5__PF1_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF1_BAR2_APERTURE_SIZE    32'h00000121
`define PCIE40E5__PF1_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_BAR2_CONTROL    32'h00000122
`define PCIE40E5__PF1_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF1_BAR3_APERTURE_SIZE    32'h00000123
`define PCIE40E5__PF1_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_BAR3_CONTROL    32'h00000124
`define PCIE40E5__PF1_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF1_BAR4_APERTURE_SIZE    32'h00000125
`define PCIE40E5__PF1_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_BAR4_CONTROL    32'h00000126
`define PCIE40E5__PF1_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF1_BAR5_APERTURE_SIZE    32'h00000127
`define PCIE40E5__PF1_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_BAR5_CONTROL    32'h00000128
`define PCIE40E5__PF1_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF1_CAPABILITY_POINTER    32'h00000129
`define PCIE40E5__PF1_CAPABILITY_POINTER_SZ 8

`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_ID    32'h0000012a
`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_ID_SZ 16

`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_LENGTH    32'h0000012b
`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_LENGTH_SZ 12

`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_NEXTPTR    32'h0000012c
`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_REVISION    32'h0000012d
`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_REVISION_SZ 4

`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_VENDOR_ID    32'h0000012e
`define PCIE40E5__PF1_CCIX_PDVSEC_CAP_VENDOR_ID_SZ 16

`define PCIE40E5__PF1_CCIX_PDVSEC_PCR_SIZE    32'h0000012f
`define PCIE40E5__PF1_CCIX_PDVSEC_PCR_SIZE_SZ 12

`define PCIE40E5__PF1_CCIX_PDVSEC_PCR_START_ADDR    32'h00000130
`define PCIE40E5__PF1_CCIX_PDVSEC_PCR_START_ADDR_SZ 12

`define PCIE40E5__PF1_CCIX_PDVSEC_PCSR_SIZE    32'h00000131
`define PCIE40E5__PF1_CCIX_PDVSEC_PCSR_SIZE_SZ 12

`define PCIE40E5__PF1_CCIX_PDVSEC_PCSR_START_ADDR    32'h00000132
`define PCIE40E5__PF1_CCIX_PDVSEC_PCSR_START_ADDR_SZ 12

`define PCIE40E5__PF1_CLASS_CODE    32'h00000133
`define PCIE40E5__PF1_CLASS_CODE_SZ 24

`define PCIE40E5__PF1_DEV_CAP_MAX_PAYLOAD_SIZE    32'h00000134
`define PCIE40E5__PF1_DEV_CAP_MAX_PAYLOAD_SIZE_SZ 3

`define PCIE40E5__PF1_DLL_FEATURE_CAP_NEXTPTR    32'h00000135
`define PCIE40E5__PF1_DLL_FEATURE_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_DSN_CAP_NEXTPTR    32'h00000136
`define PCIE40E5__PF1_DSN_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_EXPANSION_ROM_APERTURE_SIZE    32'h00000137
`define PCIE40E5__PF1_EXPANSION_ROM_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_EXPANSION_ROM_ENABLE    32'h00000138
`define PCIE40E5__PF1_EXPANSION_ROM_ENABLE_SZ 40

`define PCIE40E5__PF1_INTERRUPT_PIN    32'h00000139
`define PCIE40E5__PF1_INTERRUPT_PIN_SZ 3

`define PCIE40E5__PF1_MSIX_CAP_NEXTPTR    32'h0000013a
`define PCIE40E5__PF1_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF1_MSIX_CAP_PBA_BIR    32'h0000013b
`define PCIE40E5__PF1_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__PF1_MSIX_CAP_PBA_OFFSET    32'h0000013c
`define PCIE40E5__PF1_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__PF1_MSIX_CAP_TABLE_BIR    32'h0000013d
`define PCIE40E5__PF1_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__PF1_MSIX_CAP_TABLE_OFFSET    32'h0000013e
`define PCIE40E5__PF1_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__PF1_MSIX_CAP_TABLE_SIZE    32'h0000013f
`define PCIE40E5__PF1_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__PF1_MSI_CAP_MULTIMSGCAP    32'h00000140
`define PCIE40E5__PF1_MSI_CAP_MULTIMSGCAP_SZ 3

`define PCIE40E5__PF1_MSI_CAP_NEXTPTR    32'h00000141
`define PCIE40E5__PF1_MSI_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF1_MSI_CAP_PERVECMASKCAP    32'h00000142
`define PCIE40E5__PF1_MSI_CAP_PERVECMASKCAP_SZ 40

`define PCIE40E5__PF1_PASID_CAP_EXEC_PERM_SUPP    32'h00000143
`define PCIE40E5__PF1_PASID_CAP_EXEC_PERM_SUPP_SZ 1

`define PCIE40E5__PF1_PASID_CAP_MAX_PASID_WIDTH    32'h00000144
`define PCIE40E5__PF1_PASID_CAP_MAX_PASID_WIDTH_SZ 5

`define PCIE40E5__PF1_PASID_CAP_NEXTPTR    32'h00000145
`define PCIE40E5__PF1_PASID_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_PASID_CAP_PRIVIL_MODE_SUPP    32'h00000146
`define PCIE40E5__PF1_PASID_CAP_PRIVIL_MODE_SUPP_SZ 1

`define PCIE40E5__PF1_PCIE_CAP_NEXTPTR    32'h00000147
`define PCIE40E5__PF1_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF1_PM_CAP_NEXTPTR    32'h00000148
`define PCIE40E5__PF1_PM_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF1_PRI_CAP_NEXTPTR    32'h00000149
`define PCIE40E5__PF1_PRI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_PRI_CAP_ON    32'h0000014a
`define PCIE40E5__PF1_PRI_CAP_ON_SZ 40

`define PCIE40E5__PF1_PRI_OST_PR_CAPACITY    32'h0000014b
`define PCIE40E5__PF1_PRI_OST_PR_CAPACITY_SZ 32

`define PCIE40E5__PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED    32'h0000014c
`define PCIE40E5__PF1_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ 40

`define PCIE40E5__PF1_SRIOV_BAR0_APERTURE_SIZE    32'h0000014d
`define PCIE40E5__PF1_SRIOV_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_SRIOV_BAR0_CONTROL    32'h0000014e
`define PCIE40E5__PF1_SRIOV_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_BAR1_APERTURE_SIZE    32'h0000014f
`define PCIE40E5__PF1_SRIOV_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_SRIOV_BAR1_CONTROL    32'h00000150
`define PCIE40E5__PF1_SRIOV_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_BAR2_APERTURE_SIZE    32'h00000151
`define PCIE40E5__PF1_SRIOV_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_SRIOV_BAR2_CONTROL    32'h00000152
`define PCIE40E5__PF1_SRIOV_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_BAR3_APERTURE_SIZE    32'h00000153
`define PCIE40E5__PF1_SRIOV_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_SRIOV_BAR3_CONTROL    32'h00000154
`define PCIE40E5__PF1_SRIOV_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_BAR4_APERTURE_SIZE    32'h00000155
`define PCIE40E5__PF1_SRIOV_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF1_SRIOV_BAR4_CONTROL    32'h00000156
`define PCIE40E5__PF1_SRIOV_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_BAR5_APERTURE_SIZE    32'h00000157
`define PCIE40E5__PF1_SRIOV_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF1_SRIOV_BAR5_CONTROL    32'h00000158
`define PCIE40E5__PF1_SRIOV_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF1_SRIOV_CAP_INITIAL_VF    32'h00000159
`define PCIE40E5__PF1_SRIOV_CAP_INITIAL_VF_SZ 16

`define PCIE40E5__PF1_SRIOV_CAP_NEXTPTR    32'h0000015a
`define PCIE40E5__PF1_SRIOV_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_SRIOV_CAP_TOTAL_VF    32'h0000015b
`define PCIE40E5__PF1_SRIOV_CAP_TOTAL_VF_SZ 16

`define PCIE40E5__PF1_SRIOV_CAP_VER    32'h0000015c
`define PCIE40E5__PF1_SRIOV_CAP_VER_SZ 4

`define PCIE40E5__PF1_SRIOV_FIRST_VF_OFFSET    32'h0000015d
`define PCIE40E5__PF1_SRIOV_FIRST_VF_OFFSET_SZ 16

`define PCIE40E5__PF1_SRIOV_FUNC_DEP_LINK    32'h0000015e
`define PCIE40E5__PF1_SRIOV_FUNC_DEP_LINK_SZ 16

`define PCIE40E5__PF1_SRIOV_SUPPORTED_PAGE_SIZE    32'h0000015f
`define PCIE40E5__PF1_SRIOV_SUPPORTED_PAGE_SIZE_SZ 32

`define PCIE40E5__PF1_SRIOV_VF_DEVICE_ID    32'h00000160
`define PCIE40E5__PF1_SRIOV_VF_DEVICE_ID_SZ 16

`define PCIE40E5__PF1_TPHR_CAP_NEXTPTR    32'h00000161
`define PCIE40E5__PF1_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF1_TPHR_CAP_ST_MODE_SEL    32'h00000162
`define PCIE40E5__PF1_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__PF2_AER_CAP_NEXTPTR    32'h00000163
`define PCIE40E5__PF2_AER_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_ARI_CAP_NEXTPTR    32'h00000164
`define PCIE40E5__PF2_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_ARI_CAP_NEXT_FUNC    32'h00000165
`define PCIE40E5__PF2_ARI_CAP_NEXT_FUNC_SZ 8

`define PCIE40E5__PF2_ATS_CAP_INV_QUEUE_DEPTH    32'h00000166
`define PCIE40E5__PF2_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__PF2_ATS_CAP_NEXTPTR    32'h00000167
`define PCIE40E5__PF2_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_ATS_CAP_ON    32'h00000168
`define PCIE40E5__PF2_ATS_CAP_ON_SZ 40

`define PCIE40E5__PF2_BAR0_APERTURE_SIZE    32'h00000169
`define PCIE40E5__PF2_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_BAR0_CONTROL    32'h0000016a
`define PCIE40E5__PF2_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF2_BAR1_APERTURE_SIZE    32'h0000016b
`define PCIE40E5__PF2_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_BAR1_CONTROL    32'h0000016c
`define PCIE40E5__PF2_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF2_BAR2_APERTURE_SIZE    32'h0000016d
`define PCIE40E5__PF2_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_BAR2_CONTROL    32'h0000016e
`define PCIE40E5__PF2_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF2_BAR3_APERTURE_SIZE    32'h0000016f
`define PCIE40E5__PF2_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_BAR3_CONTROL    32'h00000170
`define PCIE40E5__PF2_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF2_BAR4_APERTURE_SIZE    32'h00000171
`define PCIE40E5__PF2_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_BAR4_CONTROL    32'h00000172
`define PCIE40E5__PF2_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF2_BAR5_APERTURE_SIZE    32'h00000173
`define PCIE40E5__PF2_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_BAR5_CONTROL    32'h00000174
`define PCIE40E5__PF2_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF2_CAPABILITY_POINTER    32'h00000175
`define PCIE40E5__PF2_CAPABILITY_POINTER_SZ 8

`define PCIE40E5__PF2_CLASS_CODE    32'h00000176
`define PCIE40E5__PF2_CLASS_CODE_SZ 24

`define PCIE40E5__PF2_DEV_CAP_MAX_PAYLOAD_SIZE    32'h00000177
`define PCIE40E5__PF2_DEV_CAP_MAX_PAYLOAD_SIZE_SZ 3

`define PCIE40E5__PF2_DLL_FEATURE_CAP_NEXTPTR    32'h00000178
`define PCIE40E5__PF2_DLL_FEATURE_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_DSN_CAP_NEXTPTR    32'h00000179
`define PCIE40E5__PF2_DSN_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_EXPANSION_ROM_APERTURE_SIZE    32'h0000017a
`define PCIE40E5__PF2_EXPANSION_ROM_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_EXPANSION_ROM_ENABLE    32'h0000017b
`define PCIE40E5__PF2_EXPANSION_ROM_ENABLE_SZ 40

`define PCIE40E5__PF2_INTERRUPT_PIN    32'h0000017c
`define PCIE40E5__PF2_INTERRUPT_PIN_SZ 3

`define PCIE40E5__PF2_MSIX_CAP_NEXTPTR    32'h0000017d
`define PCIE40E5__PF2_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF2_MSIX_CAP_PBA_BIR    32'h0000017e
`define PCIE40E5__PF2_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__PF2_MSIX_CAP_PBA_OFFSET    32'h0000017f
`define PCIE40E5__PF2_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__PF2_MSIX_CAP_TABLE_BIR    32'h00000180
`define PCIE40E5__PF2_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__PF2_MSIX_CAP_TABLE_OFFSET    32'h00000181
`define PCIE40E5__PF2_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__PF2_MSIX_CAP_TABLE_SIZE    32'h00000182
`define PCIE40E5__PF2_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__PF2_MSI_CAP_MULTIMSGCAP    32'h00000183
`define PCIE40E5__PF2_MSI_CAP_MULTIMSGCAP_SZ 3

`define PCIE40E5__PF2_MSI_CAP_NEXTPTR    32'h00000184
`define PCIE40E5__PF2_MSI_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF2_MSI_CAP_PERVECMASKCAP    32'h00000185
`define PCIE40E5__PF2_MSI_CAP_PERVECMASKCAP_SZ 40

`define PCIE40E5__PF2_PASID_CAP_EXEC_PERM_SUPP    32'h00000186
`define PCIE40E5__PF2_PASID_CAP_EXEC_PERM_SUPP_SZ 1

`define PCIE40E5__PF2_PASID_CAP_MAX_PASID_WIDTH    32'h00000187
`define PCIE40E5__PF2_PASID_CAP_MAX_PASID_WIDTH_SZ 5

`define PCIE40E5__PF2_PASID_CAP_NEXTPTR    32'h00000188
`define PCIE40E5__PF2_PASID_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_PASID_CAP_PRIVIL_MODE_SUPP    32'h00000189
`define PCIE40E5__PF2_PASID_CAP_PRIVIL_MODE_SUPP_SZ 1

`define PCIE40E5__PF2_PCIE_CAP_NEXTPTR    32'h0000018a
`define PCIE40E5__PF2_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF2_PM_CAP_NEXTPTR    32'h0000018b
`define PCIE40E5__PF2_PM_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF2_PRI_CAP_NEXTPTR    32'h0000018c
`define PCIE40E5__PF2_PRI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_PRI_CAP_ON    32'h0000018d
`define PCIE40E5__PF2_PRI_CAP_ON_SZ 40

`define PCIE40E5__PF2_PRI_OST_PR_CAPACITY    32'h0000018e
`define PCIE40E5__PF2_PRI_OST_PR_CAPACITY_SZ 32

`define PCIE40E5__PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED    32'h0000018f
`define PCIE40E5__PF2_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ 40

`define PCIE40E5__PF2_SRIOV_BAR0_APERTURE_SIZE    32'h00000190
`define PCIE40E5__PF2_SRIOV_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_SRIOV_BAR0_CONTROL    32'h00000191
`define PCIE40E5__PF2_SRIOV_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_BAR1_APERTURE_SIZE    32'h00000192
`define PCIE40E5__PF2_SRIOV_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_SRIOV_BAR1_CONTROL    32'h00000193
`define PCIE40E5__PF2_SRIOV_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_BAR2_APERTURE_SIZE    32'h00000194
`define PCIE40E5__PF2_SRIOV_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_SRIOV_BAR2_CONTROL    32'h00000195
`define PCIE40E5__PF2_SRIOV_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_BAR3_APERTURE_SIZE    32'h00000196
`define PCIE40E5__PF2_SRIOV_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_SRIOV_BAR3_CONTROL    32'h00000197
`define PCIE40E5__PF2_SRIOV_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_BAR4_APERTURE_SIZE    32'h00000198
`define PCIE40E5__PF2_SRIOV_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF2_SRIOV_BAR4_CONTROL    32'h00000199
`define PCIE40E5__PF2_SRIOV_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_BAR5_APERTURE_SIZE    32'h0000019a
`define PCIE40E5__PF2_SRIOV_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF2_SRIOV_BAR5_CONTROL    32'h0000019b
`define PCIE40E5__PF2_SRIOV_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF2_SRIOV_CAP_INITIAL_VF    32'h0000019c
`define PCIE40E5__PF2_SRIOV_CAP_INITIAL_VF_SZ 16

`define PCIE40E5__PF2_SRIOV_CAP_NEXTPTR    32'h0000019d
`define PCIE40E5__PF2_SRIOV_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_SRIOV_CAP_TOTAL_VF    32'h0000019e
`define PCIE40E5__PF2_SRIOV_CAP_TOTAL_VF_SZ 16

`define PCIE40E5__PF2_SRIOV_CAP_VER    32'h0000019f
`define PCIE40E5__PF2_SRIOV_CAP_VER_SZ 4

`define PCIE40E5__PF2_SRIOV_FIRST_VF_OFFSET    32'h000001a0
`define PCIE40E5__PF2_SRIOV_FIRST_VF_OFFSET_SZ 16

`define PCIE40E5__PF2_SRIOV_FUNC_DEP_LINK    32'h000001a1
`define PCIE40E5__PF2_SRIOV_FUNC_DEP_LINK_SZ 16

`define PCIE40E5__PF2_SRIOV_SUPPORTED_PAGE_SIZE    32'h000001a2
`define PCIE40E5__PF2_SRIOV_SUPPORTED_PAGE_SIZE_SZ 32

`define PCIE40E5__PF2_SRIOV_VF_DEVICE_ID    32'h000001a3
`define PCIE40E5__PF2_SRIOV_VF_DEVICE_ID_SZ 16

`define PCIE40E5__PF2_TPHR_CAP_NEXTPTR    32'h000001a4
`define PCIE40E5__PF2_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF2_TPHR_CAP_ST_MODE_SEL    32'h000001a5
`define PCIE40E5__PF2_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__PF3_AER_CAP_NEXTPTR    32'h000001a6
`define PCIE40E5__PF3_AER_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_ARI_CAP_NEXTPTR    32'h000001a7
`define PCIE40E5__PF3_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_ARI_CAP_NEXT_FUNC    32'h000001a8
`define PCIE40E5__PF3_ARI_CAP_NEXT_FUNC_SZ 8

`define PCIE40E5__PF3_ATS_CAP_INV_QUEUE_DEPTH    32'h000001a9
`define PCIE40E5__PF3_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__PF3_ATS_CAP_NEXTPTR    32'h000001aa
`define PCIE40E5__PF3_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_ATS_CAP_ON    32'h000001ab
`define PCIE40E5__PF3_ATS_CAP_ON_SZ 40

`define PCIE40E5__PF3_BAR0_APERTURE_SIZE    32'h000001ac
`define PCIE40E5__PF3_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_BAR0_CONTROL    32'h000001ad
`define PCIE40E5__PF3_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF3_BAR1_APERTURE_SIZE    32'h000001ae
`define PCIE40E5__PF3_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_BAR1_CONTROL    32'h000001af
`define PCIE40E5__PF3_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF3_BAR2_APERTURE_SIZE    32'h000001b0
`define PCIE40E5__PF3_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_BAR2_CONTROL    32'h000001b1
`define PCIE40E5__PF3_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF3_BAR3_APERTURE_SIZE    32'h000001b2
`define PCIE40E5__PF3_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_BAR3_CONTROL    32'h000001b3
`define PCIE40E5__PF3_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF3_BAR4_APERTURE_SIZE    32'h000001b4
`define PCIE40E5__PF3_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_BAR4_CONTROL    32'h000001b5
`define PCIE40E5__PF3_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF3_BAR5_APERTURE_SIZE    32'h000001b6
`define PCIE40E5__PF3_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_BAR5_CONTROL    32'h000001b7
`define PCIE40E5__PF3_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF3_CAPABILITY_POINTER    32'h000001b8
`define PCIE40E5__PF3_CAPABILITY_POINTER_SZ 8

`define PCIE40E5__PF3_CLASS_CODE    32'h000001b9
`define PCIE40E5__PF3_CLASS_CODE_SZ 24

`define PCIE40E5__PF3_DEV_CAP_MAX_PAYLOAD_SIZE    32'h000001ba
`define PCIE40E5__PF3_DEV_CAP_MAX_PAYLOAD_SIZE_SZ 3

`define PCIE40E5__PF3_DLL_FEATURE_CAP_NEXTPTR    32'h000001bb
`define PCIE40E5__PF3_DLL_FEATURE_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_DSN_CAP_NEXTPTR    32'h000001bc
`define PCIE40E5__PF3_DSN_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_EXPANSION_ROM_APERTURE_SIZE    32'h000001bd
`define PCIE40E5__PF3_EXPANSION_ROM_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_EXPANSION_ROM_ENABLE    32'h000001be
`define PCIE40E5__PF3_EXPANSION_ROM_ENABLE_SZ 40

`define PCIE40E5__PF3_INTERRUPT_PIN    32'h000001bf
`define PCIE40E5__PF3_INTERRUPT_PIN_SZ 3

`define PCIE40E5__PF3_MSIX_CAP_NEXTPTR    32'h000001c0
`define PCIE40E5__PF3_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF3_MSIX_CAP_PBA_BIR    32'h000001c1
`define PCIE40E5__PF3_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__PF3_MSIX_CAP_PBA_OFFSET    32'h000001c2
`define PCIE40E5__PF3_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__PF3_MSIX_CAP_TABLE_BIR    32'h000001c3
`define PCIE40E5__PF3_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__PF3_MSIX_CAP_TABLE_OFFSET    32'h000001c4
`define PCIE40E5__PF3_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__PF3_MSIX_CAP_TABLE_SIZE    32'h000001c5
`define PCIE40E5__PF3_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__PF3_MSI_CAP_MULTIMSGCAP    32'h000001c6
`define PCIE40E5__PF3_MSI_CAP_MULTIMSGCAP_SZ 3

`define PCIE40E5__PF3_MSI_CAP_NEXTPTR    32'h000001c7
`define PCIE40E5__PF3_MSI_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF3_MSI_CAP_PERVECMASKCAP    32'h000001c8
`define PCIE40E5__PF3_MSI_CAP_PERVECMASKCAP_SZ 40

`define PCIE40E5__PF3_PASID_CAP_EXEC_PERM_SUPP    32'h000001c9
`define PCIE40E5__PF3_PASID_CAP_EXEC_PERM_SUPP_SZ 1

`define PCIE40E5__PF3_PASID_CAP_MAX_PASID_WIDTH    32'h000001ca
`define PCIE40E5__PF3_PASID_CAP_MAX_PASID_WIDTH_SZ 5

`define PCIE40E5__PF3_PASID_CAP_NEXTPTR    32'h000001cb
`define PCIE40E5__PF3_PASID_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_PASID_CAP_PRIVIL_MODE_SUPP    32'h000001cc
`define PCIE40E5__PF3_PASID_CAP_PRIVIL_MODE_SUPP_SZ 1

`define PCIE40E5__PF3_PCIE_CAP_NEXTPTR    32'h000001cd
`define PCIE40E5__PF3_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF3_PM_CAP_NEXTPTR    32'h000001ce
`define PCIE40E5__PF3_PM_CAP_NEXTPTR_SZ 8

`define PCIE40E5__PF3_PRI_CAP_NEXTPTR    32'h000001cf
`define PCIE40E5__PF3_PRI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_PRI_CAP_ON    32'h000001d0
`define PCIE40E5__PF3_PRI_CAP_ON_SZ 40

`define PCIE40E5__PF3_PRI_OST_PR_CAPACITY    32'h000001d1
`define PCIE40E5__PF3_PRI_OST_PR_CAPACITY_SZ 32

`define PCIE40E5__PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED    32'h000001d2
`define PCIE40E5__PF3_SRIOV_ARI_CAPBL_HIER_PRESERVED_SZ 40

`define PCIE40E5__PF3_SRIOV_BAR0_APERTURE_SIZE    32'h000001d3
`define PCIE40E5__PF3_SRIOV_BAR0_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_SRIOV_BAR0_CONTROL    32'h000001d4
`define PCIE40E5__PF3_SRIOV_BAR0_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_BAR1_APERTURE_SIZE    32'h000001d5
`define PCIE40E5__PF3_SRIOV_BAR1_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_SRIOV_BAR1_CONTROL    32'h000001d6
`define PCIE40E5__PF3_SRIOV_BAR1_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_BAR2_APERTURE_SIZE    32'h000001d7
`define PCIE40E5__PF3_SRIOV_BAR2_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_SRIOV_BAR2_CONTROL    32'h000001d8
`define PCIE40E5__PF3_SRIOV_BAR2_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_BAR3_APERTURE_SIZE    32'h000001d9
`define PCIE40E5__PF3_SRIOV_BAR3_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_SRIOV_BAR3_CONTROL    32'h000001da
`define PCIE40E5__PF3_SRIOV_BAR3_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_BAR4_APERTURE_SIZE    32'h000001db
`define PCIE40E5__PF3_SRIOV_BAR4_APERTURE_SIZE_SZ 6

`define PCIE40E5__PF3_SRIOV_BAR4_CONTROL    32'h000001dc
`define PCIE40E5__PF3_SRIOV_BAR4_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_BAR5_APERTURE_SIZE    32'h000001dd
`define PCIE40E5__PF3_SRIOV_BAR5_APERTURE_SIZE_SZ 5

`define PCIE40E5__PF3_SRIOV_BAR5_CONTROL    32'h000001de
`define PCIE40E5__PF3_SRIOV_BAR5_CONTROL_SZ 3

`define PCIE40E5__PF3_SRIOV_CAP_INITIAL_VF    32'h000001df
`define PCIE40E5__PF3_SRIOV_CAP_INITIAL_VF_SZ 16

`define PCIE40E5__PF3_SRIOV_CAP_NEXTPTR    32'h000001e0
`define PCIE40E5__PF3_SRIOV_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_SRIOV_CAP_TOTAL_VF    32'h000001e1
`define PCIE40E5__PF3_SRIOV_CAP_TOTAL_VF_SZ 16

`define PCIE40E5__PF3_SRIOV_CAP_VER    32'h000001e2
`define PCIE40E5__PF3_SRIOV_CAP_VER_SZ 4

`define PCIE40E5__PF3_SRIOV_FIRST_VF_OFFSET    32'h000001e3
`define PCIE40E5__PF3_SRIOV_FIRST_VF_OFFSET_SZ 16

`define PCIE40E5__PF3_SRIOV_FUNC_DEP_LINK    32'h000001e4
`define PCIE40E5__PF3_SRIOV_FUNC_DEP_LINK_SZ 16

`define PCIE40E5__PF3_SRIOV_SUPPORTED_PAGE_SIZE    32'h000001e5
`define PCIE40E5__PF3_SRIOV_SUPPORTED_PAGE_SIZE_SZ 32

`define PCIE40E5__PF3_SRIOV_VF_DEVICE_ID    32'h000001e6
`define PCIE40E5__PF3_SRIOV_VF_DEVICE_ID_SZ 16

`define PCIE40E5__PF3_TPHR_CAP_NEXTPTR    32'h000001e7
`define PCIE40E5__PF3_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__PF3_TPHR_CAP_ST_MODE_SEL    32'h000001e8
`define PCIE40E5__PF3_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__PL_CCIX_ESM_CALIBRATION_TIMEOUT    32'h000001e9
`define PCIE40E5__PL_CCIX_ESM_CALIBRATION_TIMEOUT_SZ 3

`define PCIE40E5__PL_CCIX_ESM_EXTENDED_EQ_TIMEOUT    32'h000001ea
`define PCIE40E5__PL_CCIX_ESM_EXTENDED_EQ_TIMEOUT_SZ 3

`define PCIE40E5__PL_CFG_STATE_ROBUSTNESS_ENABLE    32'h000001eb
`define PCIE40E5__PL_CFG_STATE_ROBUSTNESS_ENABLE_SZ 40

`define PCIE40E5__PL_CTRL_SKP_GEN_ENABLE    32'h000001ec
`define PCIE40E5__PL_CTRL_SKP_GEN_ENABLE_SZ 40

`define PCIE40E5__PL_CTRL_SKP_PARITY_AND_CRC_CHECK_DISABLE    32'h000001ed
`define PCIE40E5__PL_CTRL_SKP_PARITY_AND_CRC_CHECK_DISABLE_SZ 40

`define PCIE40E5__PL_DEEMPH_SOURCE_SELECT    32'h000001ee
`define PCIE40E5__PL_DEEMPH_SOURCE_SELECT_SZ 40

`define PCIE40E5__PL_DESKEW_ON_SKIP_IN_GEN12    32'h000001ef
`define PCIE40E5__PL_DESKEW_ON_SKIP_IN_GEN12_SZ 40

`define PCIE40E5__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3    32'h000001f0
`define PCIE40E5__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_SZ 40

`define PCIE40E5__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4    32'h000001f1
`define PCIE40E5__PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN4_SZ 40

`define PCIE40E5__PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2    32'h000001f2
`define PCIE40E5__PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_SZ 40

`define PCIE40E5__PL_DISABLE_DC_BALANCE    32'h000001f3
`define PCIE40E5__PL_DISABLE_DC_BALANCE_SZ 40

`define PCIE40E5__PL_DISABLE_EI_INFER_IN_L0    32'h000001f4
`define PCIE40E5__PL_DISABLE_EI_INFER_IN_L0_SZ 40

`define PCIE40E5__PL_DISABLE_LANE_REVERSAL    32'h000001f5
`define PCIE40E5__PL_DISABLE_LANE_REVERSAL_SZ 40

`define PCIE40E5__PL_DISABLE_LFSR_UPDATE_ON_SKP    32'h000001f6
`define PCIE40E5__PL_DISABLE_LFSR_UPDATE_ON_SKP_SZ 2

`define PCIE40E5__PL_DISABLE_RETRAIN_ON_EB_ERROR    32'h000001f7
`define PCIE40E5__PL_DISABLE_RETRAIN_ON_EB_ERROR_SZ 40

`define PCIE40E5__PL_DISABLE_RETRAIN_ON_FRAMING_ERROR    32'h000001f8
`define PCIE40E5__PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_SZ 40

`define PCIE40E5__PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR    32'h000001f9
`define PCIE40E5__PL_DISABLE_RETRAIN_ON_SPECIFIC_FRAMING_ERROR_SZ 16

`define PCIE40E5__PL_DISABLE_UPCONFIG_CAPABLE    32'h000001fa
`define PCIE40E5__PL_DISABLE_UPCONFIG_CAPABLE_SZ 40

`define PCIE40E5__PL_ENABLE_CCIX_EDR    32'h000001fb
`define PCIE40E5__PL_ENABLE_CCIX_EDR_SZ 40

`define PCIE40E5__PL_ENABLE_CCIX_EDR_REACH_MODE    32'h000001fc
`define PCIE40E5__PL_ENABLE_CCIX_EDR_REACH_MODE_SZ 2

`define PCIE40E5__PL_EQ_ADAPT_DISABLE_COEFF_CHECK    32'h000001fd
`define PCIE40E5__PL_EQ_ADAPT_DISABLE_COEFF_CHECK_SZ 2

`define PCIE40E5__PL_EQ_ADAPT_DISABLE_PRESET_CHECK    32'h000001fe
`define PCIE40E5__PL_EQ_ADAPT_DISABLE_PRESET_CHECK_SZ 2

`define PCIE40E5__PL_EQ_ADAPT_ITER_COUNT    32'h000001ff
`define PCIE40E5__PL_EQ_ADAPT_ITER_COUNT_SZ 5

`define PCIE40E5__PL_EQ_ADAPT_REJECT_RETRY_COUNT    32'h00000200
`define PCIE40E5__PL_EQ_ADAPT_REJECT_RETRY_COUNT_SZ 2

`define PCIE40E5__PL_EQ_BYPASS_PHASE23    32'h00000201
`define PCIE40E5__PL_EQ_BYPASS_PHASE23_SZ 2

`define PCIE40E5__PL_EQ_DEFAULT_CCIX_EDR_TX_PRESET    32'h00000202
`define PCIE40E5__PL_EQ_DEFAULT_CCIX_EDR_TX_PRESET_SZ 16

`define PCIE40E5__PL_EQ_DEFAULT_RX_PRESET_HINT    32'h00000203
`define PCIE40E5__PL_EQ_DEFAULT_RX_PRESET_HINT_SZ 6

`define PCIE40E5__PL_EQ_DEFAULT_TX_PRESET    32'h00000204
`define PCIE40E5__PL_EQ_DEFAULT_TX_PRESET_SZ 16

`define PCIE40E5__PL_EQ_DISABLE_MISMATCH_CHECK    32'h00000205
`define PCIE40E5__PL_EQ_DISABLE_MISMATCH_CHECK_SZ 40

`define PCIE40E5__PL_EQ_FS    32'h00000206
`define PCIE40E5__PL_EQ_FS_SZ 6

`define PCIE40E5__PL_EQ_LF    32'h00000207
`define PCIE40E5__PL_EQ_LF_SZ 6

`define PCIE40E5__PL_EQ_LP_TXPRESET    32'h00000208
`define PCIE40E5__PL_EQ_LP_TXPRESET_SZ 16

`define PCIE40E5__PL_EQ_LP_TXPRESET2    32'h00000209
`define PCIE40E5__PL_EQ_LP_TXPRESET2_SZ 16

`define PCIE40E5__PL_EQ_RX_ADAPTATION_MODE    32'h0000020a
`define PCIE40E5__PL_EQ_RX_ADAPTATION_MODE_SZ 3

`define PCIE40E5__PL_EQ_RX_ADAPT_EQ_PHASE0    32'h0000020b
`define PCIE40E5__PL_EQ_RX_ADAPT_EQ_PHASE0_SZ 2

`define PCIE40E5__PL_EQ_RX_ADAPT_EQ_PHASE1    32'h0000020c
`define PCIE40E5__PL_EQ_RX_ADAPT_EQ_PHASE1_SZ 2

`define PCIE40E5__PL_EQ_RX_ADAPT_SIM_ENABLE    32'h0000020d
`define PCIE40E5__PL_EQ_RX_ADAPT_SIM_ENABLE_SZ 40

`define PCIE40E5__PL_EQ_RX_ADAPT_TIMER    32'h0000020e
`define PCIE40E5__PL_EQ_RX_ADAPT_TIMER_SZ 22

`define PCIE40E5__PL_EQ_RX_ADAPT_TIMER_SIM    32'h0000020f
`define PCIE40E5__PL_EQ_RX_ADAPT_TIMER_SIM_SZ 22

`define PCIE40E5__PL_EQ_RX_ADV_EQ_PER_DATA_RATE_ENABLE    32'h00000210
`define PCIE40E5__PL_EQ_RX_ADV_EQ_PER_DATA_RATE_ENABLE_SZ 4

`define PCIE40E5__PL_EQ_SHORT_ADAPT_PHASE    32'h00000211
`define PCIE40E5__PL_EQ_SHORT_ADAPT_PHASE_SZ 40

`define PCIE40E5__PL_EQ_TX_8G_EQ_TS2_ENABLE    32'h00000212
`define PCIE40E5__PL_EQ_TX_8G_EQ_TS2_ENABLE_SZ 40

`define PCIE40E5__PL_EQ_TX_MAINCUR_0    32'h00000213
`define PCIE40E5__PL_EQ_TX_MAINCUR_0_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_1    32'h00000214
`define PCIE40E5__PL_EQ_TX_MAINCUR_1_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_2    32'h00000215
`define PCIE40E5__PL_EQ_TX_MAINCUR_2_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_3    32'h00000216
`define PCIE40E5__PL_EQ_TX_MAINCUR_3_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_4    32'h00000217
`define PCIE40E5__PL_EQ_TX_MAINCUR_4_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_5    32'h00000218
`define PCIE40E5__PL_EQ_TX_MAINCUR_5_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_6    32'h00000219
`define PCIE40E5__PL_EQ_TX_MAINCUR_6_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_7    32'h0000021a
`define PCIE40E5__PL_EQ_TX_MAINCUR_7_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_8    32'h0000021b
`define PCIE40E5__PL_EQ_TX_MAINCUR_8_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_9    32'h0000021c
`define PCIE40E5__PL_EQ_TX_MAINCUR_9_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_A    32'h0000021d
`define PCIE40E5__PL_EQ_TX_MAINCUR_A_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_B    32'h0000021e
`define PCIE40E5__PL_EQ_TX_MAINCUR_B_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_C    32'h0000021f
`define PCIE40E5__PL_EQ_TX_MAINCUR_C_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_D    32'h00000220
`define PCIE40E5__PL_EQ_TX_MAINCUR_D_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_E    32'h00000221
`define PCIE40E5__PL_EQ_TX_MAINCUR_E_SZ 7

`define PCIE40E5__PL_EQ_TX_MAINCUR_F    32'h00000222
`define PCIE40E5__PL_EQ_TX_MAINCUR_F_SZ 7

`define PCIE40E5__PL_EQ_TX_POSTCUR_0    32'h00000223
`define PCIE40E5__PL_EQ_TX_POSTCUR_0_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_1    32'h00000224
`define PCIE40E5__PL_EQ_TX_POSTCUR_1_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_2    32'h00000225
`define PCIE40E5__PL_EQ_TX_POSTCUR_2_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_3    32'h00000226
`define PCIE40E5__PL_EQ_TX_POSTCUR_3_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_4    32'h00000227
`define PCIE40E5__PL_EQ_TX_POSTCUR_4_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_5    32'h00000228
`define PCIE40E5__PL_EQ_TX_POSTCUR_5_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_6    32'h00000229
`define PCIE40E5__PL_EQ_TX_POSTCUR_6_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_7    32'h0000022a
`define PCIE40E5__PL_EQ_TX_POSTCUR_7_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_8    32'h0000022b
`define PCIE40E5__PL_EQ_TX_POSTCUR_8_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_9    32'h0000022c
`define PCIE40E5__PL_EQ_TX_POSTCUR_9_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_A    32'h0000022d
`define PCIE40E5__PL_EQ_TX_POSTCUR_A_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_B    32'h0000022e
`define PCIE40E5__PL_EQ_TX_POSTCUR_B_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_C    32'h0000022f
`define PCIE40E5__PL_EQ_TX_POSTCUR_C_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_D    32'h00000230
`define PCIE40E5__PL_EQ_TX_POSTCUR_D_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_E    32'h00000231
`define PCIE40E5__PL_EQ_TX_POSTCUR_E_SZ 6

`define PCIE40E5__PL_EQ_TX_POSTCUR_F    32'h00000232
`define PCIE40E5__PL_EQ_TX_POSTCUR_F_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_0    32'h00000233
`define PCIE40E5__PL_EQ_TX_PRECUR_0_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_1    32'h00000234
`define PCIE40E5__PL_EQ_TX_PRECUR_1_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_2    32'h00000235
`define PCIE40E5__PL_EQ_TX_PRECUR_2_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_3    32'h00000236
`define PCIE40E5__PL_EQ_TX_PRECUR_3_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_4    32'h00000237
`define PCIE40E5__PL_EQ_TX_PRECUR_4_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_5    32'h00000238
`define PCIE40E5__PL_EQ_TX_PRECUR_5_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_6    32'h00000239
`define PCIE40E5__PL_EQ_TX_PRECUR_6_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_7    32'h0000023a
`define PCIE40E5__PL_EQ_TX_PRECUR_7_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_8    32'h0000023b
`define PCIE40E5__PL_EQ_TX_PRECUR_8_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_9    32'h0000023c
`define PCIE40E5__PL_EQ_TX_PRECUR_9_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_A    32'h0000023d
`define PCIE40E5__PL_EQ_TX_PRECUR_A_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_B    32'h0000023e
`define PCIE40E5__PL_EQ_TX_PRECUR_B_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_C    32'h0000023f
`define PCIE40E5__PL_EQ_TX_PRECUR_C_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_D    32'h00000240
`define PCIE40E5__PL_EQ_TX_PRECUR_D_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_E    32'h00000241
`define PCIE40E5__PL_EQ_TX_PRECUR_E_SZ 6

`define PCIE40E5__PL_EQ_TX_PRECUR_F    32'h00000242
`define PCIE40E5__PL_EQ_TX_PRECUR_F_SZ 6

`define PCIE40E5__PL_EXIT_LOOPBACK_ON_EI_ENTRY    32'h00000243
`define PCIE40E5__PL_EXIT_LOOPBACK_ON_EI_ENTRY_SZ 40

`define PCIE40E5__PL_INFER_EI_DISABLE_LPBK_ACTIVE    32'h00000244
`define PCIE40E5__PL_INFER_EI_DISABLE_LPBK_ACTIVE_SZ 40

`define PCIE40E5__PL_INFER_EI_DISABLE_REC_RC    32'h00000245
`define PCIE40E5__PL_INFER_EI_DISABLE_REC_RC_SZ 40

`define PCIE40E5__PL_INFER_EI_DISABLE_REC_SPD    32'h00000246
`define PCIE40E5__PL_INFER_EI_DISABLE_REC_SPD_SZ 40

`define PCIE40E5__PL_LANE0_CCIX_EDR_EQ_CONTROL    32'h00000247
`define PCIE40E5__PL_LANE0_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE0_EQ_CONTROL    32'h00000248
`define PCIE40E5__PL_LANE0_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE10_EQ_CONTROL    32'h00000249
`define PCIE40E5__PL_LANE10_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE11_EQ_CONTROL    32'h0000024a
`define PCIE40E5__PL_LANE11_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE12_EQ_CONTROL    32'h0000024b
`define PCIE40E5__PL_LANE12_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE13_EQ_CONTROL    32'h0000024c
`define PCIE40E5__PL_LANE13_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE14_EQ_CONTROL    32'h0000024d
`define PCIE40E5__PL_LANE14_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE15_EQ_CONTROL    32'h0000024e
`define PCIE40E5__PL_LANE15_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE1_CCIX_EDR_EQ_CONTROL    32'h0000024f
`define PCIE40E5__PL_LANE1_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE1_EQ_CONTROL    32'h00000250
`define PCIE40E5__PL_LANE1_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE2_CCIX_EDR_EQ_CONTROL    32'h00000251
`define PCIE40E5__PL_LANE2_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE2_EQ_CONTROL    32'h00000252
`define PCIE40E5__PL_LANE2_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE3_CCIX_EDR_EQ_CONTROL    32'h00000253
`define PCIE40E5__PL_LANE3_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE3_EQ_CONTROL    32'h00000254
`define PCIE40E5__PL_LANE3_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE4_CCIX_EDR_EQ_CONTROL    32'h00000255
`define PCIE40E5__PL_LANE4_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE4_EQ_CONTROL    32'h00000256
`define PCIE40E5__PL_LANE4_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE5_CCIX_EDR_EQ_CONTROL    32'h00000257
`define PCIE40E5__PL_LANE5_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE5_EQ_CONTROL    32'h00000258
`define PCIE40E5__PL_LANE5_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE6_CCIX_EDR_EQ_CONTROL    32'h00000259
`define PCIE40E5__PL_LANE6_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE6_EQ_CONTROL    32'h0000025a
`define PCIE40E5__PL_LANE6_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE7_CCIX_EDR_EQ_CONTROL    32'h0000025b
`define PCIE40E5__PL_LANE7_CCIX_EDR_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE7_EQ_CONTROL    32'h0000025c
`define PCIE40E5__PL_LANE7_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE8_EQ_CONTROL    32'h0000025d
`define PCIE40E5__PL_LANE8_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LANE9_EQ_CONTROL    32'h0000025e
`define PCIE40E5__PL_LANE9_EQ_CONTROL_SZ 32

`define PCIE40E5__PL_LINK_CAP_MAX_LINK_SPEED    32'h0000025f
`define PCIE40E5__PL_LINK_CAP_MAX_LINK_SPEED_SZ 4

`define PCIE40E5__PL_LINK_CAP_MAX_LINK_WIDTH    32'h00000260
`define PCIE40E5__PL_LINK_CAP_MAX_LINK_WIDTH_SZ 5

`define PCIE40E5__PL_N_FTS    32'h00000261
`define PCIE40E5__PL_N_FTS_SZ 8

`define PCIE40E5__PL_QUIESCE_GUARANTEE_DISABLE    32'h00000262
`define PCIE40E5__PL_QUIESCE_GUARANTEE_DISABLE_SZ 40

`define PCIE40E5__PL_RECALIBRATION_NEEDED_ON_ESM_RATE01_PROGRAMMING_CHANGE    32'h00000263
`define PCIE40E5__PL_RECALIBRATION_NEEDED_ON_ESM_RATE01_PROGRAMMING_CHANGE_SZ 40

`define PCIE40E5__PL_REDO_EQ_SOURCE_SELECT    32'h00000264
`define PCIE40E5__PL_REDO_EQ_SOURCE_SELECT_SZ 40

`define PCIE40E5__PL_REPORT_ALL_PHY_ERRORS    32'h00000265
`define PCIE40E5__PL_REPORT_ALL_PHY_ERRORS_SZ 8

`define PCIE40E5__PL_RETIMER_PRESENCE_DETECTION_SUPPORTED    32'h00000266
`define PCIE40E5__PL_RETIMER_PRESENCE_DETECTION_SUPPORTED_SZ 40

`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS    32'h00000267
`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_CLOBBER_TX_TS_SZ 2

`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_GEN3    32'h00000268
`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_GEN3_SZ 4

`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_GEN4    32'h00000269
`define PCIE40E5__PL_RX_ADAPT_TIMER_CLWS_GEN4_SZ 4

`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS    32'h0000026a
`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_CLOBBER_TX_TS_SZ 2

`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_GEN3    32'h0000026b
`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_GEN3_SZ 4

`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_GEN4    32'h0000026c
`define PCIE40E5__PL_RX_ADAPT_TIMER_RRL_GEN4_SZ 4

`define PCIE40E5__PL_RX_L0S_EXIT_TO_RECOVERY    32'h0000026d
`define PCIE40E5__PL_RX_L0S_EXIT_TO_RECOVERY_SZ 2

`define PCIE40E5__PL_SELF_TRAIN    32'h0000026e
`define PCIE40E5__PL_SELF_TRAIN_SZ 40

`define PCIE40E5__PL_SIM_FAST_LINK_TRAINING    32'h0000026f
`define PCIE40E5__PL_SIM_FAST_LINK_TRAINING_SZ 2

`define PCIE40E5__PL_SRIS_ENABLE    32'h00000270
`define PCIE40E5__PL_SRIS_ENABLE_SZ 40

`define PCIE40E5__PL_SRIS_SKPOS_GEN_SPD_VEC    32'h00000271
`define PCIE40E5__PL_SRIS_SKPOS_GEN_SPD_VEC_SZ 7

`define PCIE40E5__PL_SRIS_SKPOS_REC_SPD_VEC    32'h00000272
`define PCIE40E5__PL_SRIS_SKPOS_REC_SPD_VEC_SZ 7

`define PCIE40E5__PL_TWO_RETIMER_PRESENCE_DETECTION_SUPPORTED    32'h00000273
`define PCIE40E5__PL_TWO_RETIMER_PRESENCE_DETECTION_SUPPORTED_SZ 40

`define PCIE40E5__PL_UPSTREAM_FACING    32'h00000274
`define PCIE40E5__PL_UPSTREAM_FACING_SZ 40

`define PCIE40E5__PL_USER_SPARE    32'h00000275
`define PCIE40E5__PL_USER_SPARE_SZ 16

`define PCIE40E5__PL_USER_SPARE2    32'h00000276
`define PCIE40E5__PL_USER_SPARE2_SZ 16

`define PCIE40E5__PL_USER_SPARE3    32'h00000277
`define PCIE40E5__PL_USER_SPARE3_SZ 32

`define PCIE40E5__PM_ASPML0S_TIMEOUT    32'h00000278
`define PCIE40E5__PM_ASPML0S_TIMEOUT_SZ 16

`define PCIE40E5__PM_ASPML1_ENTRY_DELAY    32'h00000279
`define PCIE40E5__PM_ASPML1_ENTRY_DELAY_SZ 20

`define PCIE40E5__PM_ENABLE_L23_ENTRY    32'h0000027a
`define PCIE40E5__PM_ENABLE_L23_ENTRY_SZ 40

`define PCIE40E5__PM_ENABLE_SLOT_POWER_CAPTURE    32'h0000027b
`define PCIE40E5__PM_ENABLE_SLOT_POWER_CAPTURE_SZ 40

`define PCIE40E5__PM_L1_REENTRY_DELAY    32'h0000027c
`define PCIE40E5__PM_L1_REENTRY_DELAY_SZ 32

`define PCIE40E5__PM_PME_TURNOFF_ACK_DELAY    32'h0000027d
`define PCIE40E5__PM_PME_TURNOFF_ACK_DELAY_SZ 16

`define PCIE40E5__ROOT_CAP_CRS_SW_VISIBILITY    32'h0000027e
`define PCIE40E5__ROOT_CAP_CRS_SW_VISIBILITY_SZ 40

`define PCIE40E5__SIM_DEVICE    32'h0000027f
`define PCIE40E5__SIM_DEVICE_SZ 144

`define PCIE40E5__SPARE_BIT0    32'h00000280
`define PCIE40E5__SPARE_BIT0_SZ 40

`define PCIE40E5__SPARE_BIT1    32'h00000281
`define PCIE40E5__SPARE_BIT1_SZ 1

`define PCIE40E5__SPARE_BIT2    32'h00000282
`define PCIE40E5__SPARE_BIT2_SZ 1

`define PCIE40E5__SPARE_BIT3    32'h00000283
`define PCIE40E5__SPARE_BIT3_SZ 40

`define PCIE40E5__SPARE_BIT4    32'h00000284
`define PCIE40E5__SPARE_BIT4_SZ 1

`define PCIE40E5__SPARE_BIT5    32'h00000285
`define PCIE40E5__SPARE_BIT5_SZ 1

`define PCIE40E5__SPARE_BIT6    32'h00000286
`define PCIE40E5__SPARE_BIT6_SZ 1

`define PCIE40E5__SPARE_BIT7    32'h00000287
`define PCIE40E5__SPARE_BIT7_SZ 1

`define PCIE40E5__SPARE_BIT8    32'h00000288
`define PCIE40E5__SPARE_BIT8_SZ 1

`define PCIE40E5__SPARE_BYTE0    32'h00000289
`define PCIE40E5__SPARE_BYTE0_SZ 8

`define PCIE40E5__SPARE_BYTE1    32'h0000028a
`define PCIE40E5__SPARE_BYTE1_SZ 8

`define PCIE40E5__SPARE_BYTE2    32'h0000028b
`define PCIE40E5__SPARE_BYTE2_SZ 8

`define PCIE40E5__SPARE_BYTE3    32'h0000028c
`define PCIE40E5__SPARE_BYTE3_SZ 8

`define PCIE40E5__SPARE_WORD0    32'h0000028d
`define PCIE40E5__SPARE_WORD0_SZ 32

`define PCIE40E5__SPARE_WORD1    32'h0000028e
`define PCIE40E5__SPARE_WORD1_SZ 32

`define PCIE40E5__SPARE_WORD2    32'h0000028f
`define PCIE40E5__SPARE_WORD2_SZ 32

`define PCIE40E5__SPARE_WORD3    32'h00000290
`define PCIE40E5__SPARE_WORD3_SZ 32

`define PCIE40E5__SRIOV_CAP_ENABLE    32'h00000291
`define PCIE40E5__SRIOV_CAP_ENABLE_SZ 4

`define PCIE40E5__TL2CFG_IF_PARITY_CHK    32'h00000292
`define PCIE40E5__TL2CFG_IF_PARITY_CHK_SZ 40

`define PCIE40E5__TL_COMPLETION_RAM_NUM_TLPS    32'h00000293
`define PCIE40E5__TL_COMPLETION_RAM_NUM_TLPS_SZ 2

`define PCIE40E5__TL_COMPLETION_RAM_SIZE    32'h00000294
`define PCIE40E5__TL_COMPLETION_RAM_SIZE_SZ 2

`define PCIE40E5__TL_CREDITS_CD    32'h00000295
`define PCIE40E5__TL_CREDITS_CD_SZ 12

`define PCIE40E5__TL_CREDITS_CD_VC1    32'h00000296
`define PCIE40E5__TL_CREDITS_CD_VC1_SZ 12

`define PCIE40E5__TL_CREDITS_CH    32'h00000297
`define PCIE40E5__TL_CREDITS_CH_SZ 8

`define PCIE40E5__TL_CREDITS_CH_VC1    32'h00000298
`define PCIE40E5__TL_CREDITS_CH_VC1_SZ 8

`define PCIE40E5__TL_CREDITS_NPD    32'h00000299
`define PCIE40E5__TL_CREDITS_NPD_SZ 12

`define PCIE40E5__TL_CREDITS_NPD_VC1    32'h0000029a
`define PCIE40E5__TL_CREDITS_NPD_VC1_SZ 12

`define PCIE40E5__TL_CREDITS_NPH    32'h0000029b
`define PCIE40E5__TL_CREDITS_NPH_SZ 8

`define PCIE40E5__TL_CREDITS_NPH_VC1    32'h0000029c
`define PCIE40E5__TL_CREDITS_NPH_VC1_SZ 8

`define PCIE40E5__TL_CREDITS_PD    32'h0000029d
`define PCIE40E5__TL_CREDITS_PD_SZ 12

`define PCIE40E5__TL_CREDITS_PD_VC1    32'h0000029e
`define PCIE40E5__TL_CREDITS_PD_VC1_SZ 12

`define PCIE40E5__TL_CREDITS_PH    32'h0000029f
`define PCIE40E5__TL_CREDITS_PH_SZ 8

`define PCIE40E5__TL_CREDITS_PH_VC1    32'h000002a0
`define PCIE40E5__TL_CREDITS_PH_VC1_SZ 8

`define PCIE40E5__TL_DISABLE_RX_FLOW_CTL    32'h000002a1
`define PCIE40E5__TL_DISABLE_RX_FLOW_CTL_SZ 40

`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TIME    32'h000002a2
`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TIME_SZ 5

`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TIME_VC1    32'h000002a3
`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TIME_VC1_SZ 5

`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT    32'h000002a4
`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT_SZ 5

`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT_VC1    32'h000002a5
`define PCIE40E5__TL_FC_UPDATE_MIN_INTERVAL_TLP_COUNT_VC1_SZ 5

`define PCIE40E5__TL_FEATURE_ENABLE_FC_SCALING    32'h000002a6
`define PCIE40E5__TL_FEATURE_ENABLE_FC_SCALING_SZ 40

`define PCIE40E5__TL_NP_FIFO_NUM_TLPS    32'h000002a7
`define PCIE40E5__TL_NP_FIFO_NUM_TLPS_SZ 1

`define PCIE40E5__TL_PF_ENABLE_REG    32'h000002a8
`define PCIE40E5__TL_PF_ENABLE_REG_SZ 2

`define PCIE40E5__TL_POSTED_RAM_SIZE    32'h000002a9
`define PCIE40E5__TL_POSTED_RAM_SIZE_SZ 1

`define PCIE40E5__TL_RX_CCIX_FIFO_FROM_RAM_READ_PIPELINE    32'h000002aa
`define PCIE40E5__TL_RX_CCIX_FIFO_FROM_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_CCIX_FIFO_RAM_SIZE    32'h000002ab
`define PCIE40E5__TL_RX_CCIX_FIFO_RAM_SIZE_SZ 1

`define PCIE40E5__TL_RX_CCIX_FIFO_TO_RAM_READ_PIPELINE    32'h000002ac
`define PCIE40E5__TL_RX_CCIX_FIFO_TO_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_CCIX_FIFO_TO_RAM_WRITE_PIPELINE    32'h000002ad
`define PCIE40E5__TL_RX_CCIX_FIFO_TO_RAM_WRITE_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE    32'h000002ae
`define PCIE40E5__TL_RX_COMPLETION_FROM_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_COMPLETION_TO_RAM_READ_PIPELINE    32'h000002af
`define PCIE40E5__TL_RX_COMPLETION_TO_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE    32'h000002b0
`define PCIE40E5__TL_RX_COMPLETION_TO_RAM_WRITE_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_POSTED_FROM_RAM_READ_PIPELINE    32'h000002b1
`define PCIE40E5__TL_RX_POSTED_FROM_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_POSTED_TO_RAM_READ_PIPELINE    32'h000002b2
`define PCIE40E5__TL_RX_POSTED_TO_RAM_READ_PIPELINE_SZ 40

`define PCIE40E5__TL_RX_POSTED_TO_RAM_WRITE_PIPELINE    32'h000002b3
`define PCIE40E5__TL_RX_POSTED_TO_RAM_WRITE_PIPELINE_SZ 40

`define PCIE40E5__TL_TX_MUX_STRICT_PRIORITY    32'h000002b4
`define PCIE40E5__TL_TX_MUX_STRICT_PRIORITY_SZ 40

`define PCIE40E5__TL_TX_TLP_STRADDLE_ENABLE    32'h000002b5
`define PCIE40E5__TL_TX_TLP_STRADDLE_ENABLE_SZ 40

`define PCIE40E5__TL_TX_TLP_TERMINATE_PARITY    32'h000002b6
`define PCIE40E5__TL_TX_TLP_TERMINATE_PARITY_SZ 40

`define PCIE40E5__TL_USER_SPARE    32'h000002b7
`define PCIE40E5__TL_USER_SPARE_SZ 16

`define PCIE40E5__TPH_FROM_RAM_PIPELINE    32'h000002b8
`define PCIE40E5__TPH_FROM_RAM_PIPELINE_SZ 40

`define PCIE40E5__TPH_TO_RAM_PIPELINE    32'h000002b9
`define PCIE40E5__TPH_TO_RAM_PIPELINE_SZ 40

`define PCIE40E5__VC1_BASE_DISABLE    32'h000002ba
`define PCIE40E5__VC1_BASE_DISABLE_SZ 40

`define PCIE40E5__VF0_CAPABILITY_POINTER    32'h000002bb
`define PCIE40E5__VF0_CAPABILITY_POINTER_SZ 8

`define PCIE40E5__VFG0_10B_TAG_REQUESTER_SUPPORTED    32'h000002bc
`define PCIE40E5__VFG0_10B_TAG_REQUESTER_SUPPORTED_SZ 40

`define PCIE40E5__VFG0_ARI_CAP_NEXTPTR    32'h000002bd
`define PCIE40E5__VFG0_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG0_ATS_CAP_INV_QUEUE_DEPTH    32'h000002be
`define PCIE40E5__VFG0_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__VFG0_ATS_CAP_NEXTPTR    32'h000002bf
`define PCIE40E5__VFG0_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG0_ATS_CAP_ON    32'h000002c0
`define PCIE40E5__VFG0_ATS_CAP_ON_SZ 40

`define PCIE40E5__VFG0_MSIX_CAP_NEXTPTR    32'h000002c1
`define PCIE40E5__VFG0_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG0_MSIX_CAP_PBA_BIR    32'h000002c2
`define PCIE40E5__VFG0_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__VFG0_MSIX_CAP_PBA_OFFSET    32'h000002c3
`define PCIE40E5__VFG0_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__VFG0_MSIX_CAP_TABLE_BIR    32'h000002c4
`define PCIE40E5__VFG0_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__VFG0_MSIX_CAP_TABLE_OFFSET    32'h000002c5
`define PCIE40E5__VFG0_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__VFG0_MSIX_CAP_TABLE_SIZE    32'h000002c6
`define PCIE40E5__VFG0_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__VFG0_PCIE_CAP_NEXTPTR    32'h000002c7
`define PCIE40E5__VFG0_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG0_TPHR_CAP_NEXTPTR    32'h000002c8
`define PCIE40E5__VFG0_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG0_TPHR_CAP_ST_MODE_SEL    32'h000002c9
`define PCIE40E5__VFG0_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__VFG1_10B_TAG_REQUESTER_SUPPORTED    32'h000002ca
`define PCIE40E5__VFG1_10B_TAG_REQUESTER_SUPPORTED_SZ 40

`define PCIE40E5__VFG1_ARI_CAP_NEXTPTR    32'h000002cb
`define PCIE40E5__VFG1_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG1_ATS_CAP_INV_QUEUE_DEPTH    32'h000002cc
`define PCIE40E5__VFG1_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__VFG1_ATS_CAP_NEXTPTR    32'h000002cd
`define PCIE40E5__VFG1_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG1_ATS_CAP_ON    32'h000002ce
`define PCIE40E5__VFG1_ATS_CAP_ON_SZ 40

`define PCIE40E5__VFG1_MSIX_CAP_NEXTPTR    32'h000002cf
`define PCIE40E5__VFG1_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG1_MSIX_CAP_PBA_BIR    32'h000002d0
`define PCIE40E5__VFG1_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__VFG1_MSIX_CAP_PBA_OFFSET    32'h000002d1
`define PCIE40E5__VFG1_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__VFG1_MSIX_CAP_TABLE_BIR    32'h000002d2
`define PCIE40E5__VFG1_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__VFG1_MSIX_CAP_TABLE_OFFSET    32'h000002d3
`define PCIE40E5__VFG1_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__VFG1_MSIX_CAP_TABLE_SIZE    32'h000002d4
`define PCIE40E5__VFG1_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__VFG1_PCIE_CAP_NEXTPTR    32'h000002d5
`define PCIE40E5__VFG1_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG1_TPHR_CAP_NEXTPTR    32'h000002d6
`define PCIE40E5__VFG1_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG1_TPHR_CAP_ST_MODE_SEL    32'h000002d7
`define PCIE40E5__VFG1_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__VFG2_10B_TAG_REQUESTER_SUPPORTED    32'h000002d8
`define PCIE40E5__VFG2_10B_TAG_REQUESTER_SUPPORTED_SZ 40

`define PCIE40E5__VFG2_ARI_CAP_NEXTPTR    32'h000002d9
`define PCIE40E5__VFG2_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG2_ATS_CAP_INV_QUEUE_DEPTH    32'h000002da
`define PCIE40E5__VFG2_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__VFG2_ATS_CAP_NEXTPTR    32'h000002db
`define PCIE40E5__VFG2_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG2_ATS_CAP_ON    32'h000002dc
`define PCIE40E5__VFG2_ATS_CAP_ON_SZ 40

`define PCIE40E5__VFG2_MSIX_CAP_NEXTPTR    32'h000002dd
`define PCIE40E5__VFG2_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG2_MSIX_CAP_PBA_BIR    32'h000002de
`define PCIE40E5__VFG2_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__VFG2_MSIX_CAP_PBA_OFFSET    32'h000002df
`define PCIE40E5__VFG2_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__VFG2_MSIX_CAP_TABLE_BIR    32'h000002e0
`define PCIE40E5__VFG2_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__VFG2_MSIX_CAP_TABLE_OFFSET    32'h000002e1
`define PCIE40E5__VFG2_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__VFG2_MSIX_CAP_TABLE_SIZE    32'h000002e2
`define PCIE40E5__VFG2_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__VFG2_PCIE_CAP_NEXTPTR    32'h000002e3
`define PCIE40E5__VFG2_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG2_TPHR_CAP_NEXTPTR    32'h000002e4
`define PCIE40E5__VFG2_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG2_TPHR_CAP_ST_MODE_SEL    32'h000002e5
`define PCIE40E5__VFG2_TPHR_CAP_ST_MODE_SEL_SZ 3

`define PCIE40E5__VFG3_10B_TAG_REQUESTER_SUPPORTED    32'h000002e6
`define PCIE40E5__VFG3_10B_TAG_REQUESTER_SUPPORTED_SZ 40

`define PCIE40E5__VFG3_ARI_CAP_NEXTPTR    32'h000002e7
`define PCIE40E5__VFG3_ARI_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG3_ATS_CAP_INV_QUEUE_DEPTH    32'h000002e8
`define PCIE40E5__VFG3_ATS_CAP_INV_QUEUE_DEPTH_SZ 5

`define PCIE40E5__VFG3_ATS_CAP_NEXTPTR    32'h000002e9
`define PCIE40E5__VFG3_ATS_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG3_ATS_CAP_ON    32'h000002ea
`define PCIE40E5__VFG3_ATS_CAP_ON_SZ 40

`define PCIE40E5__VFG3_MSIX_CAP_NEXTPTR    32'h000002eb
`define PCIE40E5__VFG3_MSIX_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG3_MSIX_CAP_PBA_BIR    32'h000002ec
`define PCIE40E5__VFG3_MSIX_CAP_PBA_BIR_SZ 3

`define PCIE40E5__VFG3_MSIX_CAP_PBA_OFFSET    32'h000002ed
`define PCIE40E5__VFG3_MSIX_CAP_PBA_OFFSET_SZ 29

`define PCIE40E5__VFG3_MSIX_CAP_TABLE_BIR    32'h000002ee
`define PCIE40E5__VFG3_MSIX_CAP_TABLE_BIR_SZ 3

`define PCIE40E5__VFG3_MSIX_CAP_TABLE_OFFSET    32'h000002ef
`define PCIE40E5__VFG3_MSIX_CAP_TABLE_OFFSET_SZ 29

`define PCIE40E5__VFG3_MSIX_CAP_TABLE_SIZE    32'h000002f0
`define PCIE40E5__VFG3_MSIX_CAP_TABLE_SIZE_SZ 11

`define PCIE40E5__VFG3_PCIE_CAP_NEXTPTR    32'h000002f1
`define PCIE40E5__VFG3_PCIE_CAP_NEXTPTR_SZ 8

`define PCIE40E5__VFG3_TPHR_CAP_NEXTPTR    32'h000002f2
`define PCIE40E5__VFG3_TPHR_CAP_NEXTPTR_SZ 12

`define PCIE40E5__VFG3_TPHR_CAP_ST_MODE_SEL    32'h000002f3
`define PCIE40E5__VFG3_TPHR_CAP_ST_MODE_SEL_SZ 3

`endif  // B_PCIE40E5_DEFINES_VH