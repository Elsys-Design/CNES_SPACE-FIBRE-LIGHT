`include "B_DSP_OUTPUT58_defines.vh"

reg [`DSP_OUTPUT58_DATA_SZ-1:0] ATTR [0:`DSP_OUTPUT58_ADDR_N-1];
reg [`DSP_OUTPUT58__ADREG_SZ-1:0] ADREG_REG = ADREG;
reg [`DSP_OUTPUT58__AMULTSEL_SZ:1] AMULTSEL_REG = AMULTSEL;
reg [`DSP_OUTPUT58__AUTORESET_PATDET_SZ:1] AUTORESET_PATDET_REG = AUTORESET_PATDET;
reg [`DSP_OUTPUT58__AUTORESET_PRIORITY_SZ:1] AUTORESET_PRIORITY_REG = AUTORESET_PRIORITY;
reg [`DSP_OUTPUT58__BMULTSEL_SZ:1] BMULTSEL_REG = BMULTSEL;
reg [`DSP_OUTPUT58__DSP_MODE_SZ:1] DSP_MODE_REG = DSP_MODE;
reg IS_RSTP_INVERTED_REG = IS_RSTP_INVERTED;
reg [`DSP_OUTPUT58__LEGACY_SZ:1] LEGACY_REG = LEGACY;
reg [`DSP_OUTPUT58__PREG_SZ-1:0] PREG_REG = PREG;
reg [`DSP_OUTPUT58__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;
reg [`DSP_OUTPUT58__USE_MULT_SZ:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_OUTPUT58__ADREG] = ADREG;
  ATTR[`DSP_OUTPUT58__AMULTSEL] = AMULTSEL;
  ATTR[`DSP_OUTPUT58__AUTORESET_PATDET] = AUTORESET_PATDET;
  ATTR[`DSP_OUTPUT58__AUTORESET_PRIORITY] = AUTORESET_PRIORITY;
  ATTR[`DSP_OUTPUT58__BMULTSEL] = BMULTSEL;
  ATTR[`DSP_OUTPUT58__DSP_MODE] = DSP_MODE;
  ATTR[`DSP_OUTPUT58__IS_RSTP_INVERTED] = IS_RSTP_INVERTED;
  ATTR[`DSP_OUTPUT58__LEGACY] = LEGACY;
  ATTR[`DSP_OUTPUT58__PREG] = PREG;
  ATTR[`DSP_OUTPUT58__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_OUTPUT58__USE_MULT] = USE_MULT;
end

always @(*) begin
  ADREG_REG = ATTR[`DSP_OUTPUT58__ADREG];
  AMULTSEL_REG = ATTR[`DSP_OUTPUT58__AMULTSEL];
  AUTORESET_PATDET_REG = ATTR[`DSP_OUTPUT58__AUTORESET_PATDET];
  AUTORESET_PRIORITY_REG = ATTR[`DSP_OUTPUT58__AUTORESET_PRIORITY];
  BMULTSEL_REG = ATTR[`DSP_OUTPUT58__BMULTSEL];
  DSP_MODE_REG = ATTR[`DSP_OUTPUT58__DSP_MODE];
  IS_RSTP_INVERTED_REG = ATTR[`DSP_OUTPUT58__IS_RSTP_INVERTED];
  LEGACY_REG = ATTR[`DSP_OUTPUT58__LEGACY];
  PREG_REG = ATTR[`DSP_OUTPUT58__PREG];
  RESET_MODE_REG = ATTR[`DSP_OUTPUT58__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_OUTPUT58__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_OUTPUT58_ADDR_SZ-1:0] addr;
  input  [`DSP_OUTPUT58_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_OUTPUT58_DATA_SZ-1:0] read_attr;
  input  [`DSP_OUTPUT58_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
