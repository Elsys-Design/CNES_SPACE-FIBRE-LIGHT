// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_URAM288_DEFINES_VH
`else
`define B_URAM288_DEFINES_VH

// Look-up table parameters
//

`define URAM288_ADDR_N  38
`define URAM288_ADDR_SZ 32
`define URAM288_DATA_SZ 144

// Attribute addresses
//

`define URAM288__AUTO_SLEEP_LATENCY    32'h00000000
`define URAM288__AUTO_SLEEP_LATENCY_SZ 32

`define URAM288__AVG_CONS_INACTIVE_CYCLES    32'h00000001
`define URAM288__AVG_CONS_INACTIVE_CYCLES_SZ 32

`define URAM288__BWE_MODE_A    32'h00000002
`define URAM288__BWE_MODE_A_SZ 144

`define URAM288__BWE_MODE_B    32'h00000003
`define URAM288__BWE_MODE_B_SZ 144

`define URAM288__CASCADE_ORDER_A    32'h00000004
`define URAM288__CASCADE_ORDER_A_SZ 48

`define URAM288__CASCADE_ORDER_B    32'h00000005
`define URAM288__CASCADE_ORDER_B_SZ 48

`define URAM288__EN_AUTO_SLEEP_MODE    32'h00000006
`define URAM288__EN_AUTO_SLEEP_MODE_SZ 40

`define URAM288__EN_ECC_RD_A    32'h00000007
`define URAM288__EN_ECC_RD_A_SZ 40

`define URAM288__EN_ECC_RD_B    32'h00000008
`define URAM288__EN_ECC_RD_B_SZ 40

`define URAM288__EN_ECC_WR_A    32'h00000009
`define URAM288__EN_ECC_WR_A_SZ 40

`define URAM288__EN_ECC_WR_B    32'h0000000a
`define URAM288__EN_ECC_WR_B_SZ 40

`define URAM288__IREG_PRE_A    32'h0000000b
`define URAM288__IREG_PRE_A_SZ 40

`define URAM288__IREG_PRE_B    32'h0000000c
`define URAM288__IREG_PRE_B_SZ 40

`define URAM288__IS_CLK_INVERTED    32'h0000000d
`define URAM288__IS_CLK_INVERTED_SZ 1

`define URAM288__IS_EN_A_INVERTED    32'h0000000e
`define URAM288__IS_EN_A_INVERTED_SZ 1

`define URAM288__IS_EN_B_INVERTED    32'h0000000f
`define URAM288__IS_EN_B_INVERTED_SZ 1

`define URAM288__IS_RDB_WR_A_INVERTED    32'h00000010
`define URAM288__IS_RDB_WR_A_INVERTED_SZ 1

`define URAM288__IS_RDB_WR_B_INVERTED    32'h00000011
`define URAM288__IS_RDB_WR_B_INVERTED_SZ 1

`define URAM288__IS_RST_A_INVERTED    32'h00000012
`define URAM288__IS_RST_A_INVERTED_SZ 1

`define URAM288__IS_RST_B_INVERTED    32'h00000013
`define URAM288__IS_RST_B_INVERTED_SZ 1

`define URAM288__MATRIX_ID    32'h00000014
`define URAM288__MATRIX_ID_SZ 32

`define URAM288__NUM_UNIQUE_SELF_ADDR_A    32'h00000015
`define URAM288__NUM_UNIQUE_SELF_ADDR_A_SZ 32

`define URAM288__NUM_UNIQUE_SELF_ADDR_B    32'h00000016
`define URAM288__NUM_UNIQUE_SELF_ADDR_B_SZ 32

`define URAM288__NUM_URAM_IN_MATRIX    32'h00000017
`define URAM288__NUM_URAM_IN_MATRIX_SZ 32

`define URAM288__OREG_A    32'h00000018
`define URAM288__OREG_A_SZ 40

`define URAM288__OREG_B    32'h00000019
`define URAM288__OREG_B_SZ 40

`define URAM288__OREG_ECC_A    32'h0000001a
`define URAM288__OREG_ECC_A_SZ 40

`define URAM288__OREG_ECC_B    32'h0000001b
`define URAM288__OREG_ECC_B_SZ 40

`define URAM288__REG_CAS_A    32'h0000001c
`define URAM288__REG_CAS_A_SZ 40

`define URAM288__REG_CAS_B    32'h0000001d
`define URAM288__REG_CAS_B_SZ 40

`define URAM288__RST_MODE_A    32'h0000001e
`define URAM288__RST_MODE_A_SZ 40

`define URAM288__RST_MODE_B    32'h0000001f
`define URAM288__RST_MODE_B_SZ 40

`define URAM288__SELF_ADDR_A    32'h00000020
`define URAM288__SELF_ADDR_A_SZ 11

`define URAM288__SELF_ADDR_B    32'h00000021
`define URAM288__SELF_ADDR_B_SZ 11

`define URAM288__SELF_MASK_A    32'h00000022
`define URAM288__SELF_MASK_A_SZ 11

`define URAM288__SELF_MASK_B    32'h00000023
`define URAM288__SELF_MASK_B_SZ 11

`define URAM288__USE_EXT_CE_A    32'h00000024
`define URAM288__USE_EXT_CE_A_SZ 40

`define URAM288__USE_EXT_CE_B    32'h00000025
`define URAM288__USE_EXT_CE_B_SZ 40

`endif  // B_URAM288_DEFINES_VH