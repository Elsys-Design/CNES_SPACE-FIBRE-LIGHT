// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_A_B_DATA58_DEFINES_VH
`else
`define B_DSP_A_B_DATA58_DEFINES_VH

// Look-up table parameters
//

`define DSP_A_B_DATA58_ADDR_N  12
`define DSP_A_B_DATA58_ADDR_SZ 32
`define DSP_A_B_DATA58_DATA_SZ 56

// Attribute addresses
//

`define DSP_A_B_DATA58__ACASCREG    32'h00000000
`define DSP_A_B_DATA58__ACASCREG_SZ 32

`define DSP_A_B_DATA58__AMULTSEL    32'h00000001
`define DSP_A_B_DATA58__AMULTSEL_SZ 16

`define DSP_A_B_DATA58__AREG    32'h00000002
`define DSP_A_B_DATA58__AREG_SZ 32

`define DSP_A_B_DATA58__A_INPUT    32'h00000003
`define DSP_A_B_DATA58__A_INPUT_SZ 56

`define DSP_A_B_DATA58__BCASCREG    32'h00000004
`define DSP_A_B_DATA58__BCASCREG_SZ 32

`define DSP_A_B_DATA58__BMULTSEL    32'h00000005
`define DSP_A_B_DATA58__BMULTSEL_SZ 16

`define DSP_A_B_DATA58__BREG    32'h00000006
`define DSP_A_B_DATA58__BREG_SZ 32

`define DSP_A_B_DATA58__B_INPUT    32'h00000007
`define DSP_A_B_DATA58__B_INPUT_SZ 56

`define DSP_A_B_DATA58__DSP_MODE    32'h00000008
`define DSP_A_B_DATA58__DSP_MODE_SZ 48

`define DSP_A_B_DATA58__IS_RSTA_INVERTED    32'h00000009
`define DSP_A_B_DATA58__IS_RSTA_INVERTED_SZ 1

`define DSP_A_B_DATA58__IS_RSTB_INVERTED    32'h0000000a
`define DSP_A_B_DATA58__IS_RSTB_INVERTED_SZ 1

`define DSP_A_B_DATA58__RESET_MODE    32'h0000000b
`define DSP_A_B_DATA58__RESET_MODE_SZ 40

`endif  // B_DSP_A_B_DATA58_DEFINES_VH