`include "B_NOC_NCRB_defines.vh"

reg [`NOC_NCRB_DATA_SZ-1:0] ATTR [0:`NOC_NCRB_ADDR_N-1];
reg [`NOC_NCRB__REG_P0_0_VCA_TOKEN_SZ-1:0] REG_P0_0_VCA_TOKEN_REG = REG_P0_0_VCA_TOKEN;
reg [`NOC_NCRB__REG_P0_1_VCA_TOKEN_SZ-1:0] REG_P0_1_VCA_TOKEN_REG = REG_P0_1_VCA_TOKEN;
reg [`NOC_NCRB__REG_P0_R2W_EB_CTRL_SZ-1:0] REG_P0_R2W_EB_CTRL_REG = REG_P0_R2W_EB_CTRL;
reg [`NOC_NCRB__REG_P0_W2R_EB_CTRL_SZ-1:0] REG_P0_W2R_EB_CTRL_REG = REG_P0_W2R_EB_CTRL;
reg [`NOC_NCRB__REG_P1_0_VCA_TOKEN_SZ-1:0] REG_P1_0_VCA_TOKEN_REG = REG_P1_0_VCA_TOKEN;
reg [`NOC_NCRB__REG_P1_1_VCA_TOKEN_SZ-1:0] REG_P1_1_VCA_TOKEN_REG = REG_P1_1_VCA_TOKEN;
reg [`NOC_NCRB__REG_P1_R2W_EB_CTRL_SZ-1:0] REG_P1_R2W_EB_CTRL_REG = REG_P1_R2W_EB_CTRL;
reg [`NOC_NCRB__REG_P1_W2R_EB_CTRL_SZ-1:0] REG_P1_W2R_EB_CTRL_REG = REG_P1_W2R_EB_CTRL;
reg REG_PIPE_MODE_REG = REG_PIPE_MODE;

initial begin
  ATTR[`NOC_NCRB__REG_P0_0_VCA_TOKEN] = REG_P0_0_VCA_TOKEN;
  ATTR[`NOC_NCRB__REG_P0_1_VCA_TOKEN] = REG_P0_1_VCA_TOKEN;
  ATTR[`NOC_NCRB__REG_P0_R2W_EB_CTRL] = REG_P0_R2W_EB_CTRL;
  ATTR[`NOC_NCRB__REG_P0_W2R_EB_CTRL] = REG_P0_W2R_EB_CTRL;
  ATTR[`NOC_NCRB__REG_P1_0_VCA_TOKEN] = REG_P1_0_VCA_TOKEN;
  ATTR[`NOC_NCRB__REG_P1_1_VCA_TOKEN] = REG_P1_1_VCA_TOKEN;
  ATTR[`NOC_NCRB__REG_P1_R2W_EB_CTRL] = REG_P1_R2W_EB_CTRL;
  ATTR[`NOC_NCRB__REG_P1_W2R_EB_CTRL] = REG_P1_W2R_EB_CTRL;
  ATTR[`NOC_NCRB__REG_PIPE_MODE] = REG_PIPE_MODE;
end

always @(trig_attr) begin
  REG_P0_0_VCA_TOKEN_REG = ATTR[`NOC_NCRB__REG_P0_0_VCA_TOKEN];
  REG_P0_1_VCA_TOKEN_REG = ATTR[`NOC_NCRB__REG_P0_1_VCA_TOKEN];
  REG_P0_R2W_EB_CTRL_REG = ATTR[`NOC_NCRB__REG_P0_R2W_EB_CTRL];
  REG_P0_W2R_EB_CTRL_REG = ATTR[`NOC_NCRB__REG_P0_W2R_EB_CTRL];
  REG_P1_0_VCA_TOKEN_REG = ATTR[`NOC_NCRB__REG_P1_0_VCA_TOKEN];
  REG_P1_1_VCA_TOKEN_REG = ATTR[`NOC_NCRB__REG_P1_1_VCA_TOKEN];
  REG_P1_R2W_EB_CTRL_REG = ATTR[`NOC_NCRB__REG_P1_R2W_EB_CTRL];
  REG_P1_W2R_EB_CTRL_REG = ATTR[`NOC_NCRB__REG_P1_W2R_EB_CTRL];
  REG_PIPE_MODE_REG = ATTR[`NOC_NCRB__REG_PIPE_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`NOC_NCRB_ADDR_SZ-1:0] addr;
  input  [`NOC_NCRB_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`NOC_NCRB_DATA_SZ-1:0] read_attr;
  input  [`NOC_NCRB_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
