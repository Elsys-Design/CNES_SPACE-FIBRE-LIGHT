// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DDRMC_DEFINES_VH
`else
`define B_DDRMC_DEFINES_VH

// Look-up table parameters
//

`define DDRMC_ADDR_N  782
`define DDRMC_ADDR_SZ 32
`define DDRMC_DATA_SZ 144

// Attribute addresses
//

`define DDRMC__ARBITER_CONFIG    32'h00000000
`define DDRMC__ARBITER_CONFIG_SZ 1

`define DDRMC__CAL_CS_CH    32'h00000001
`define DDRMC__CAL_CS_CH_SZ 2

`define DDRMC__CAL_MODE    32'h00000002
`define DDRMC__CAL_MODE_SZ 1

`define DDRMC__CHANNELS    32'h00000003
`define DDRMC__CHANNELS_SZ 32

`define DDRMC__CLK_GATE    32'h00000004
`define DDRMC__CLK_GATE_SZ 19

`define DDRMC__COMMAND_BUS_OPTION    32'h00000005
`define DDRMC__COMMAND_BUS_OPTION_SZ 144

`define DDRMC__CPLX_BURST_ARRAY0    32'h00000006
`define DDRMC__CPLX_BURST_ARRAY0_SZ 5

`define DDRMC__CPLX_BURST_ARRAY1    32'h00000007
`define DDRMC__CPLX_BURST_ARRAY1_SZ 5

`define DDRMC__CPLX_BURST_ARRAY10    32'h00000008
`define DDRMC__CPLX_BURST_ARRAY10_SZ 5

`define DDRMC__CPLX_BURST_ARRAY11    32'h00000009
`define DDRMC__CPLX_BURST_ARRAY11_SZ 5

`define DDRMC__CPLX_BURST_ARRAY12    32'h0000000a
`define DDRMC__CPLX_BURST_ARRAY12_SZ 5

`define DDRMC__CPLX_BURST_ARRAY13    32'h0000000b
`define DDRMC__CPLX_BURST_ARRAY13_SZ 5

`define DDRMC__CPLX_BURST_ARRAY14    32'h0000000c
`define DDRMC__CPLX_BURST_ARRAY14_SZ 5

`define DDRMC__CPLX_BURST_ARRAY15    32'h0000000d
`define DDRMC__CPLX_BURST_ARRAY15_SZ 5

`define DDRMC__CPLX_BURST_ARRAY16    32'h0000000e
`define DDRMC__CPLX_BURST_ARRAY16_SZ 5

`define DDRMC__CPLX_BURST_ARRAY17    32'h0000000f
`define DDRMC__CPLX_BURST_ARRAY17_SZ 5

`define DDRMC__CPLX_BURST_ARRAY18    32'h00000010
`define DDRMC__CPLX_BURST_ARRAY18_SZ 5

`define DDRMC__CPLX_BURST_ARRAY19    32'h00000011
`define DDRMC__CPLX_BURST_ARRAY19_SZ 5

`define DDRMC__CPLX_BURST_ARRAY2    32'h00000012
`define DDRMC__CPLX_BURST_ARRAY2_SZ 5

`define DDRMC__CPLX_BURST_ARRAY20    32'h00000013
`define DDRMC__CPLX_BURST_ARRAY20_SZ 5

`define DDRMC__CPLX_BURST_ARRAY21    32'h00000014
`define DDRMC__CPLX_BURST_ARRAY21_SZ 5

`define DDRMC__CPLX_BURST_ARRAY22    32'h00000015
`define DDRMC__CPLX_BURST_ARRAY22_SZ 5

`define DDRMC__CPLX_BURST_ARRAY3    32'h00000016
`define DDRMC__CPLX_BURST_ARRAY3_SZ 5

`define DDRMC__CPLX_BURST_ARRAY4    32'h00000017
`define DDRMC__CPLX_BURST_ARRAY4_SZ 5

`define DDRMC__CPLX_BURST_ARRAY5    32'h00000018
`define DDRMC__CPLX_BURST_ARRAY5_SZ 5

`define DDRMC__CPLX_BURST_ARRAY6    32'h00000019
`define DDRMC__CPLX_BURST_ARRAY6_SZ 5

`define DDRMC__CPLX_BURST_ARRAY7    32'h0000001a
`define DDRMC__CPLX_BURST_ARRAY7_SZ 5

`define DDRMC__CPLX_BURST_ARRAY8    32'h0000001b
`define DDRMC__CPLX_BURST_ARRAY8_SZ 5

`define DDRMC__CPLX_BURST_ARRAY9    32'h0000001c
`define DDRMC__CPLX_BURST_ARRAY9_SZ 5

`define DDRMC__CPLX_CONFIG    32'h0000001d
`define DDRMC__CPLX_CONFIG_SZ 31

`define DDRMC__CPLX_CONFIG2    32'h0000001e
`define DDRMC__CPLX_CONFIG2_SZ 25

`define DDRMC__CPLX_CONFIG3    32'h0000001f
`define DDRMC__CPLX_CONFIG3_SZ 10

`define DDRMC__CPLX_PATTERN0    32'h00000020
`define DDRMC__CPLX_PATTERN0_SZ 16

`define DDRMC__CPLX_PATTERN1    32'h00000021
`define DDRMC__CPLX_PATTERN1_SZ 16

`define DDRMC__CPLX_PATTERN10    32'h00000022
`define DDRMC__CPLX_PATTERN10_SZ 16

`define DDRMC__CPLX_PATTERN100    32'h00000023
`define DDRMC__CPLX_PATTERN100_SZ 16

`define DDRMC__CPLX_PATTERN101    32'h00000024
`define DDRMC__CPLX_PATTERN101_SZ 16

`define DDRMC__CPLX_PATTERN102    32'h00000025
`define DDRMC__CPLX_PATTERN102_SZ 16

`define DDRMC__CPLX_PATTERN103    32'h00000026
`define DDRMC__CPLX_PATTERN103_SZ 16

`define DDRMC__CPLX_PATTERN104    32'h00000027
`define DDRMC__CPLX_PATTERN104_SZ 16

`define DDRMC__CPLX_PATTERN105    32'h00000028
`define DDRMC__CPLX_PATTERN105_SZ 16

`define DDRMC__CPLX_PATTERN106    32'h00000029
`define DDRMC__CPLX_PATTERN106_SZ 16

`define DDRMC__CPLX_PATTERN107    32'h0000002a
`define DDRMC__CPLX_PATTERN107_SZ 16

`define DDRMC__CPLX_PATTERN108    32'h0000002b
`define DDRMC__CPLX_PATTERN108_SZ 16

`define DDRMC__CPLX_PATTERN109    32'h0000002c
`define DDRMC__CPLX_PATTERN109_SZ 16

`define DDRMC__CPLX_PATTERN11    32'h0000002d
`define DDRMC__CPLX_PATTERN11_SZ 16

`define DDRMC__CPLX_PATTERN110    32'h0000002e
`define DDRMC__CPLX_PATTERN110_SZ 16

`define DDRMC__CPLX_PATTERN111    32'h0000002f
`define DDRMC__CPLX_PATTERN111_SZ 16

`define DDRMC__CPLX_PATTERN112    32'h00000030
`define DDRMC__CPLX_PATTERN112_SZ 16

`define DDRMC__CPLX_PATTERN113    32'h00000031
`define DDRMC__CPLX_PATTERN113_SZ 16

`define DDRMC__CPLX_PATTERN114    32'h00000032
`define DDRMC__CPLX_PATTERN114_SZ 16

`define DDRMC__CPLX_PATTERN115    32'h00000033
`define DDRMC__CPLX_PATTERN115_SZ 16

`define DDRMC__CPLX_PATTERN116    32'h00000034
`define DDRMC__CPLX_PATTERN116_SZ 16

`define DDRMC__CPLX_PATTERN117    32'h00000035
`define DDRMC__CPLX_PATTERN117_SZ 16

`define DDRMC__CPLX_PATTERN118    32'h00000036
`define DDRMC__CPLX_PATTERN118_SZ 16

`define DDRMC__CPLX_PATTERN119    32'h00000037
`define DDRMC__CPLX_PATTERN119_SZ 16

`define DDRMC__CPLX_PATTERN12    32'h00000038
`define DDRMC__CPLX_PATTERN12_SZ 16

`define DDRMC__CPLX_PATTERN120    32'h00000039
`define DDRMC__CPLX_PATTERN120_SZ 16

`define DDRMC__CPLX_PATTERN121    32'h0000003a
`define DDRMC__CPLX_PATTERN121_SZ 16

`define DDRMC__CPLX_PATTERN122    32'h0000003b
`define DDRMC__CPLX_PATTERN122_SZ 16

`define DDRMC__CPLX_PATTERN123    32'h0000003c
`define DDRMC__CPLX_PATTERN123_SZ 16

`define DDRMC__CPLX_PATTERN124    32'h0000003d
`define DDRMC__CPLX_PATTERN124_SZ 16

`define DDRMC__CPLX_PATTERN125    32'h0000003e
`define DDRMC__CPLX_PATTERN125_SZ 16

`define DDRMC__CPLX_PATTERN126    32'h0000003f
`define DDRMC__CPLX_PATTERN126_SZ 16

`define DDRMC__CPLX_PATTERN127    32'h00000040
`define DDRMC__CPLX_PATTERN127_SZ 16

`define DDRMC__CPLX_PATTERN128    32'h00000041
`define DDRMC__CPLX_PATTERN128_SZ 16

`define DDRMC__CPLX_PATTERN129    32'h00000042
`define DDRMC__CPLX_PATTERN129_SZ 16

`define DDRMC__CPLX_PATTERN13    32'h00000043
`define DDRMC__CPLX_PATTERN13_SZ 16

`define DDRMC__CPLX_PATTERN130    32'h00000044
`define DDRMC__CPLX_PATTERN130_SZ 16

`define DDRMC__CPLX_PATTERN131    32'h00000045
`define DDRMC__CPLX_PATTERN131_SZ 16

`define DDRMC__CPLX_PATTERN132    32'h00000046
`define DDRMC__CPLX_PATTERN132_SZ 16

`define DDRMC__CPLX_PATTERN133    32'h00000047
`define DDRMC__CPLX_PATTERN133_SZ 16

`define DDRMC__CPLX_PATTERN134    32'h00000048
`define DDRMC__CPLX_PATTERN134_SZ 16

`define DDRMC__CPLX_PATTERN135    32'h00000049
`define DDRMC__CPLX_PATTERN135_SZ 16

`define DDRMC__CPLX_PATTERN136    32'h0000004a
`define DDRMC__CPLX_PATTERN136_SZ 16

`define DDRMC__CPLX_PATTERN137    32'h0000004b
`define DDRMC__CPLX_PATTERN137_SZ 16

`define DDRMC__CPLX_PATTERN138    32'h0000004c
`define DDRMC__CPLX_PATTERN138_SZ 16

`define DDRMC__CPLX_PATTERN139    32'h0000004d
`define DDRMC__CPLX_PATTERN139_SZ 16

`define DDRMC__CPLX_PATTERN14    32'h0000004e
`define DDRMC__CPLX_PATTERN14_SZ 16

`define DDRMC__CPLX_PATTERN140    32'h0000004f
`define DDRMC__CPLX_PATTERN140_SZ 16

`define DDRMC__CPLX_PATTERN141    32'h00000050
`define DDRMC__CPLX_PATTERN141_SZ 16

`define DDRMC__CPLX_PATTERN142    32'h00000051
`define DDRMC__CPLX_PATTERN142_SZ 16

`define DDRMC__CPLX_PATTERN143    32'h00000052
`define DDRMC__CPLX_PATTERN143_SZ 16

`define DDRMC__CPLX_PATTERN144    32'h00000053
`define DDRMC__CPLX_PATTERN144_SZ 16

`define DDRMC__CPLX_PATTERN145    32'h00000054
`define DDRMC__CPLX_PATTERN145_SZ 16

`define DDRMC__CPLX_PATTERN146    32'h00000055
`define DDRMC__CPLX_PATTERN146_SZ 16

`define DDRMC__CPLX_PATTERN147    32'h00000056
`define DDRMC__CPLX_PATTERN147_SZ 16

`define DDRMC__CPLX_PATTERN148    32'h00000057
`define DDRMC__CPLX_PATTERN148_SZ 16

`define DDRMC__CPLX_PATTERN149    32'h00000058
`define DDRMC__CPLX_PATTERN149_SZ 16

`define DDRMC__CPLX_PATTERN15    32'h00000059
`define DDRMC__CPLX_PATTERN15_SZ 16

`define DDRMC__CPLX_PATTERN150    32'h0000005a
`define DDRMC__CPLX_PATTERN150_SZ 16

`define DDRMC__CPLX_PATTERN151    32'h0000005b
`define DDRMC__CPLX_PATTERN151_SZ 16

`define DDRMC__CPLX_PATTERN152    32'h0000005c
`define DDRMC__CPLX_PATTERN152_SZ 16

`define DDRMC__CPLX_PATTERN153    32'h0000005d
`define DDRMC__CPLX_PATTERN153_SZ 16

`define DDRMC__CPLX_PATTERN154    32'h0000005e
`define DDRMC__CPLX_PATTERN154_SZ 16

`define DDRMC__CPLX_PATTERN155    32'h0000005f
`define DDRMC__CPLX_PATTERN155_SZ 16

`define DDRMC__CPLX_PATTERN156    32'h00000060
`define DDRMC__CPLX_PATTERN156_SZ 16

`define DDRMC__CPLX_PATTERN16    32'h00000061
`define DDRMC__CPLX_PATTERN16_SZ 16

`define DDRMC__CPLX_PATTERN17    32'h00000062
`define DDRMC__CPLX_PATTERN17_SZ 16

`define DDRMC__CPLX_PATTERN18    32'h00000063
`define DDRMC__CPLX_PATTERN18_SZ 16

`define DDRMC__CPLX_PATTERN19    32'h00000064
`define DDRMC__CPLX_PATTERN19_SZ 16

`define DDRMC__CPLX_PATTERN2    32'h00000065
`define DDRMC__CPLX_PATTERN2_SZ 16

`define DDRMC__CPLX_PATTERN20    32'h00000066
`define DDRMC__CPLX_PATTERN20_SZ 16

`define DDRMC__CPLX_PATTERN21    32'h00000067
`define DDRMC__CPLX_PATTERN21_SZ 16

`define DDRMC__CPLX_PATTERN22    32'h00000068
`define DDRMC__CPLX_PATTERN22_SZ 16

`define DDRMC__CPLX_PATTERN23    32'h00000069
`define DDRMC__CPLX_PATTERN23_SZ 16

`define DDRMC__CPLX_PATTERN24    32'h0000006a
`define DDRMC__CPLX_PATTERN24_SZ 16

`define DDRMC__CPLX_PATTERN25    32'h0000006b
`define DDRMC__CPLX_PATTERN25_SZ 16

`define DDRMC__CPLX_PATTERN26    32'h0000006c
`define DDRMC__CPLX_PATTERN26_SZ 16

`define DDRMC__CPLX_PATTERN27    32'h0000006d
`define DDRMC__CPLX_PATTERN27_SZ 16

`define DDRMC__CPLX_PATTERN28    32'h0000006e
`define DDRMC__CPLX_PATTERN28_SZ 16

`define DDRMC__CPLX_PATTERN29    32'h0000006f
`define DDRMC__CPLX_PATTERN29_SZ 16

`define DDRMC__CPLX_PATTERN3    32'h00000070
`define DDRMC__CPLX_PATTERN3_SZ 16

`define DDRMC__CPLX_PATTERN30    32'h00000071
`define DDRMC__CPLX_PATTERN30_SZ 16

`define DDRMC__CPLX_PATTERN31    32'h00000072
`define DDRMC__CPLX_PATTERN31_SZ 16

`define DDRMC__CPLX_PATTERN32    32'h00000073
`define DDRMC__CPLX_PATTERN32_SZ 16

`define DDRMC__CPLX_PATTERN33    32'h00000074
`define DDRMC__CPLX_PATTERN33_SZ 16

`define DDRMC__CPLX_PATTERN34    32'h00000075
`define DDRMC__CPLX_PATTERN34_SZ 16

`define DDRMC__CPLX_PATTERN35    32'h00000076
`define DDRMC__CPLX_PATTERN35_SZ 16

`define DDRMC__CPLX_PATTERN36    32'h00000077
`define DDRMC__CPLX_PATTERN36_SZ 16

`define DDRMC__CPLX_PATTERN37    32'h00000078
`define DDRMC__CPLX_PATTERN37_SZ 16

`define DDRMC__CPLX_PATTERN38    32'h00000079
`define DDRMC__CPLX_PATTERN38_SZ 16

`define DDRMC__CPLX_PATTERN39    32'h0000007a
`define DDRMC__CPLX_PATTERN39_SZ 16

`define DDRMC__CPLX_PATTERN4    32'h0000007b
`define DDRMC__CPLX_PATTERN4_SZ 16

`define DDRMC__CPLX_PATTERN40    32'h0000007c
`define DDRMC__CPLX_PATTERN40_SZ 16

`define DDRMC__CPLX_PATTERN41    32'h0000007d
`define DDRMC__CPLX_PATTERN41_SZ 16

`define DDRMC__CPLX_PATTERN42    32'h0000007e
`define DDRMC__CPLX_PATTERN42_SZ 16

`define DDRMC__CPLX_PATTERN43    32'h0000007f
`define DDRMC__CPLX_PATTERN43_SZ 16

`define DDRMC__CPLX_PATTERN44    32'h00000080
`define DDRMC__CPLX_PATTERN44_SZ 16

`define DDRMC__CPLX_PATTERN45    32'h00000081
`define DDRMC__CPLX_PATTERN45_SZ 16

`define DDRMC__CPLX_PATTERN46    32'h00000082
`define DDRMC__CPLX_PATTERN46_SZ 16

`define DDRMC__CPLX_PATTERN47    32'h00000083
`define DDRMC__CPLX_PATTERN47_SZ 16

`define DDRMC__CPLX_PATTERN48    32'h00000084
`define DDRMC__CPLX_PATTERN48_SZ 16

`define DDRMC__CPLX_PATTERN49    32'h00000085
`define DDRMC__CPLX_PATTERN49_SZ 16

`define DDRMC__CPLX_PATTERN5    32'h00000086
`define DDRMC__CPLX_PATTERN5_SZ 16

`define DDRMC__CPLX_PATTERN50    32'h00000087
`define DDRMC__CPLX_PATTERN50_SZ 16

`define DDRMC__CPLX_PATTERN51    32'h00000088
`define DDRMC__CPLX_PATTERN51_SZ 16

`define DDRMC__CPLX_PATTERN52    32'h00000089
`define DDRMC__CPLX_PATTERN52_SZ 16

`define DDRMC__CPLX_PATTERN53    32'h0000008a
`define DDRMC__CPLX_PATTERN53_SZ 16

`define DDRMC__CPLX_PATTERN54    32'h0000008b
`define DDRMC__CPLX_PATTERN54_SZ 16

`define DDRMC__CPLX_PATTERN55    32'h0000008c
`define DDRMC__CPLX_PATTERN55_SZ 16

`define DDRMC__CPLX_PATTERN56    32'h0000008d
`define DDRMC__CPLX_PATTERN56_SZ 16

`define DDRMC__CPLX_PATTERN57    32'h0000008e
`define DDRMC__CPLX_PATTERN57_SZ 16

`define DDRMC__CPLX_PATTERN58    32'h0000008f
`define DDRMC__CPLX_PATTERN58_SZ 16

`define DDRMC__CPLX_PATTERN59    32'h00000090
`define DDRMC__CPLX_PATTERN59_SZ 16

`define DDRMC__CPLX_PATTERN6    32'h00000091
`define DDRMC__CPLX_PATTERN6_SZ 16

`define DDRMC__CPLX_PATTERN60    32'h00000092
`define DDRMC__CPLX_PATTERN60_SZ 16

`define DDRMC__CPLX_PATTERN61    32'h00000093
`define DDRMC__CPLX_PATTERN61_SZ 16

`define DDRMC__CPLX_PATTERN62    32'h00000094
`define DDRMC__CPLX_PATTERN62_SZ 16

`define DDRMC__CPLX_PATTERN63    32'h00000095
`define DDRMC__CPLX_PATTERN63_SZ 16

`define DDRMC__CPLX_PATTERN64    32'h00000096
`define DDRMC__CPLX_PATTERN64_SZ 16

`define DDRMC__CPLX_PATTERN65    32'h00000097
`define DDRMC__CPLX_PATTERN65_SZ 16

`define DDRMC__CPLX_PATTERN66    32'h00000098
`define DDRMC__CPLX_PATTERN66_SZ 16

`define DDRMC__CPLX_PATTERN67    32'h00000099
`define DDRMC__CPLX_PATTERN67_SZ 16

`define DDRMC__CPLX_PATTERN68    32'h0000009a
`define DDRMC__CPLX_PATTERN68_SZ 16

`define DDRMC__CPLX_PATTERN69    32'h0000009b
`define DDRMC__CPLX_PATTERN69_SZ 16

`define DDRMC__CPLX_PATTERN7    32'h0000009c
`define DDRMC__CPLX_PATTERN7_SZ 16

`define DDRMC__CPLX_PATTERN70    32'h0000009d
`define DDRMC__CPLX_PATTERN70_SZ 16

`define DDRMC__CPLX_PATTERN71    32'h0000009e
`define DDRMC__CPLX_PATTERN71_SZ 16

`define DDRMC__CPLX_PATTERN72    32'h0000009f
`define DDRMC__CPLX_PATTERN72_SZ 16

`define DDRMC__CPLX_PATTERN73    32'h000000a0
`define DDRMC__CPLX_PATTERN73_SZ 16

`define DDRMC__CPLX_PATTERN74    32'h000000a1
`define DDRMC__CPLX_PATTERN74_SZ 16

`define DDRMC__CPLX_PATTERN75    32'h000000a2
`define DDRMC__CPLX_PATTERN75_SZ 16

`define DDRMC__CPLX_PATTERN76    32'h000000a3
`define DDRMC__CPLX_PATTERN76_SZ 16

`define DDRMC__CPLX_PATTERN77    32'h000000a4
`define DDRMC__CPLX_PATTERN77_SZ 16

`define DDRMC__CPLX_PATTERN78    32'h000000a5
`define DDRMC__CPLX_PATTERN78_SZ 16

`define DDRMC__CPLX_PATTERN79    32'h000000a6
`define DDRMC__CPLX_PATTERN79_SZ 16

`define DDRMC__CPLX_PATTERN8    32'h000000a7
`define DDRMC__CPLX_PATTERN8_SZ 16

`define DDRMC__CPLX_PATTERN80    32'h000000a8
`define DDRMC__CPLX_PATTERN80_SZ 16

`define DDRMC__CPLX_PATTERN81    32'h000000a9
`define DDRMC__CPLX_PATTERN81_SZ 16

`define DDRMC__CPLX_PATTERN82    32'h000000aa
`define DDRMC__CPLX_PATTERN82_SZ 16

`define DDRMC__CPLX_PATTERN83    32'h000000ab
`define DDRMC__CPLX_PATTERN83_SZ 16

`define DDRMC__CPLX_PATTERN84    32'h000000ac
`define DDRMC__CPLX_PATTERN84_SZ 16

`define DDRMC__CPLX_PATTERN85    32'h000000ad
`define DDRMC__CPLX_PATTERN85_SZ 16

`define DDRMC__CPLX_PATTERN86    32'h000000ae
`define DDRMC__CPLX_PATTERN86_SZ 16

`define DDRMC__CPLX_PATTERN87    32'h000000af
`define DDRMC__CPLX_PATTERN87_SZ 16

`define DDRMC__CPLX_PATTERN88    32'h000000b0
`define DDRMC__CPLX_PATTERN88_SZ 16

`define DDRMC__CPLX_PATTERN89    32'h000000b1
`define DDRMC__CPLX_PATTERN89_SZ 16

`define DDRMC__CPLX_PATTERN9    32'h000000b2
`define DDRMC__CPLX_PATTERN9_SZ 16

`define DDRMC__CPLX_PATTERN90    32'h000000b3
`define DDRMC__CPLX_PATTERN90_SZ 16

`define DDRMC__CPLX_PATTERN91    32'h000000b4
`define DDRMC__CPLX_PATTERN91_SZ 16

`define DDRMC__CPLX_PATTERN92    32'h000000b5
`define DDRMC__CPLX_PATTERN92_SZ 16

`define DDRMC__CPLX_PATTERN93    32'h000000b6
`define DDRMC__CPLX_PATTERN93_SZ 16

`define DDRMC__CPLX_PATTERN94    32'h000000b7
`define DDRMC__CPLX_PATTERN94_SZ 16

`define DDRMC__CPLX_PATTERN95    32'h000000b8
`define DDRMC__CPLX_PATTERN95_SZ 16

`define DDRMC__CPLX_PATTERN96    32'h000000b9
`define DDRMC__CPLX_PATTERN96_SZ 16

`define DDRMC__CPLX_PATTERN97    32'h000000ba
`define DDRMC__CPLX_PATTERN97_SZ 16

`define DDRMC__CPLX_PATTERN98    32'h000000bb
`define DDRMC__CPLX_PATTERN98_SZ 16

`define DDRMC__CPLX_PATTERN99    32'h000000bc
`define DDRMC__CPLX_PATTERN99_SZ 16

`define DDRMC__DATA_RATE    32'h000000bd
`define DDRMC__DATA_RATE_SZ 64

`define DDRMC__DATA_WIDTH    32'h000000be
`define DDRMC__DATA_WIDTH_SZ 32

`define DDRMC__DBG_TRIGGER    32'h000000bf
`define DDRMC__DBG_TRIGGER_SZ 3

`define DDRMC__DC_CMD_CREDITS    32'h000000c0
`define DDRMC__DC_CMD_CREDITS_SZ 12

`define DDRMC__DDR_MODE    32'h000000c1
`define DDRMC__DDR_MODE_SZ 48

`define DDRMC__DEFAULT_PATTERN    32'h000000c2
`define DDRMC__DEFAULT_PATTERN_SZ 10

`define DDRMC__ECC_USAGE    32'h000000c3
`define DDRMC__ECC_USAGE_SZ 40

`define DDRMC__EXMON_CLR_EXE    32'h000000c4
`define DDRMC__EXMON_CLR_EXE_SZ 9

`define DDRMC__FIFO_RDEN    32'h000000c5
`define DDRMC__FIFO_RDEN_SZ 7

`define DDRMC__INPUT_TERMINATION    32'h000000c6
`define DDRMC__INPUT_TERMINATION_SZ 32

`define DDRMC__OUTPUT_TERMINATION    32'h000000c7
`define DDRMC__OUTPUT_TERMINATION_SZ 32

`define DDRMC__PHY_RANK_READ_OVERRIDE    32'h000000c8
`define DDRMC__PHY_RANK_READ_OVERRIDE_SZ 18

`define DDRMC__PHY_RANK_WRITE_OVERRIDE    32'h000000c9
`define DDRMC__PHY_RANK_WRITE_OVERRIDE_SZ 18

`define DDRMC__PHY_RDEN0    32'h000000ca
`define DDRMC__PHY_RDEN0_SZ 7

`define DDRMC__PHY_RDEN1    32'h000000cb
`define DDRMC__PHY_RDEN1_SZ 7

`define DDRMC__PHY_RDEN10    32'h000000cc
`define DDRMC__PHY_RDEN10_SZ 7

`define DDRMC__PHY_RDEN11    32'h000000cd
`define DDRMC__PHY_RDEN11_SZ 7

`define DDRMC__PHY_RDEN12    32'h000000ce
`define DDRMC__PHY_RDEN12_SZ 7

`define DDRMC__PHY_RDEN13    32'h000000cf
`define DDRMC__PHY_RDEN13_SZ 7

`define DDRMC__PHY_RDEN14    32'h000000d0
`define DDRMC__PHY_RDEN14_SZ 7

`define DDRMC__PHY_RDEN15    32'h000000d1
`define DDRMC__PHY_RDEN15_SZ 7

`define DDRMC__PHY_RDEN16    32'h000000d2
`define DDRMC__PHY_RDEN16_SZ 7

`define DDRMC__PHY_RDEN17    32'h000000d3
`define DDRMC__PHY_RDEN17_SZ 7

`define DDRMC__PHY_RDEN18    32'h000000d4
`define DDRMC__PHY_RDEN18_SZ 7

`define DDRMC__PHY_RDEN19    32'h000000d5
`define DDRMC__PHY_RDEN19_SZ 7

`define DDRMC__PHY_RDEN2    32'h000000d6
`define DDRMC__PHY_RDEN2_SZ 7

`define DDRMC__PHY_RDEN20    32'h000000d7
`define DDRMC__PHY_RDEN20_SZ 7

`define DDRMC__PHY_RDEN21    32'h000000d8
`define DDRMC__PHY_RDEN21_SZ 7

`define DDRMC__PHY_RDEN22    32'h000000d9
`define DDRMC__PHY_RDEN22_SZ 7

`define DDRMC__PHY_RDEN23    32'h000000da
`define DDRMC__PHY_RDEN23_SZ 7

`define DDRMC__PHY_RDEN24    32'h000000db
`define DDRMC__PHY_RDEN24_SZ 7

`define DDRMC__PHY_RDEN25    32'h000000dc
`define DDRMC__PHY_RDEN25_SZ 7

`define DDRMC__PHY_RDEN26    32'h000000dd
`define DDRMC__PHY_RDEN26_SZ 7

`define DDRMC__PHY_RDEN3    32'h000000de
`define DDRMC__PHY_RDEN3_SZ 7

`define DDRMC__PHY_RDEN4    32'h000000df
`define DDRMC__PHY_RDEN4_SZ 7

`define DDRMC__PHY_RDEN5    32'h000000e0
`define DDRMC__PHY_RDEN5_SZ 7

`define DDRMC__PHY_RDEN6    32'h000000e1
`define DDRMC__PHY_RDEN6_SZ 7

`define DDRMC__PHY_RDEN7    32'h000000e2
`define DDRMC__PHY_RDEN7_SZ 7

`define DDRMC__PHY_RDEN8    32'h000000e3
`define DDRMC__PHY_RDEN8_SZ 7

`define DDRMC__PHY_RDEN9    32'h000000e4
`define DDRMC__PHY_RDEN9_SZ 7

`define DDRMC__PRBS_CNT    32'h000000e5
`define DDRMC__PRBS_CNT_SZ 32

`define DDRMC__PRBS_CONFIG    32'h000000e6
`define DDRMC__PRBS_CONFIG_SZ 17

`define DDRMC__PRBS_CONFIG2    32'h000000e7
`define DDRMC__PRBS_CONFIG2_SZ 18

`define DDRMC__PRBS_SEED0    32'h000000e8
`define DDRMC__PRBS_SEED0_SZ 23

`define DDRMC__PRBS_SEED1    32'h000000e9
`define DDRMC__PRBS_SEED1_SZ 23

`define DDRMC__PRBS_SEED2    32'h000000ea
`define DDRMC__PRBS_SEED2_SZ 23

`define DDRMC__PRBS_SEED3    32'h000000eb
`define DDRMC__PRBS_SEED3_SZ 23

`define DDRMC__PRBS_SEED4    32'h000000ec
`define DDRMC__PRBS_SEED4_SZ 23

`define DDRMC__PRBS_SEED5    32'h000000ed
`define DDRMC__PRBS_SEED5_SZ 23

`define DDRMC__PRBS_SEED6    32'h000000ee
`define DDRMC__PRBS_SEED6_SZ 23

`define DDRMC__PRBS_SEED7    32'h000000ef
`define DDRMC__PRBS_SEED7_SZ 23

`define DDRMC__PRBS_SEED8    32'h000000f0
`define DDRMC__PRBS_SEED8_SZ 23

`define DDRMC__RAM_SETTING_RF2PHS    32'h000000f1
`define DDRMC__RAM_SETTING_RF2PHS_SZ 8

`define DDRMC__RAM_SETTING_RFSPHD    32'h000000f2
`define DDRMC__RAM_SETTING_RFSPHD_SZ 7

`define DDRMC__RAM_SETTING_SRSPHD    32'h000000f3
`define DDRMC__RAM_SETTING_SRSPHD_SZ 7

`define DDRMC__READ_BANDWIDTH    32'h000000f4
`define DDRMC__READ_BANDWIDTH_SZ 64

`define DDRMC__REG_ADEC0    32'h000000f5
`define DDRMC__REG_ADEC0_SZ 20

`define DDRMC__REG_ADEC1    32'h000000f6
`define DDRMC__REG_ADEC1_SZ 20

`define DDRMC__REG_ADEC10    32'h000000f7
`define DDRMC__REG_ADEC10_SZ 30

`define DDRMC__REG_ADEC11    32'h000000f8
`define DDRMC__REG_ADEC11_SZ 24

`define DDRMC__REG_ADEC2    32'h000000f9
`define DDRMC__REG_ADEC2_SZ 21

`define DDRMC__REG_ADEC3    32'h000000fa
`define DDRMC__REG_ADEC3_SZ 20

`define DDRMC__REG_ADEC4    32'h000000fb
`define DDRMC__REG_ADEC4_SZ 30

`define DDRMC__REG_ADEC5    32'h000000fc
`define DDRMC__REG_ADEC5_SZ 30

`define DDRMC__REG_ADEC6    32'h000000fd
`define DDRMC__REG_ADEC6_SZ 30

`define DDRMC__REG_ADEC7    32'h000000fe
`define DDRMC__REG_ADEC7_SZ 30

`define DDRMC__REG_ADEC8    32'h000000ff
`define DDRMC__REG_ADEC8_SZ 30

`define DDRMC__REG_ADEC9    32'h00000100
`define DDRMC__REG_ADEC9_SZ 30

`define DDRMC__REG_CMDQ_BER_RATE_CTRL    32'h00000101
`define DDRMC__REG_CMDQ_BER_RATE_CTRL_SZ 22

`define DDRMC__REG_CMDQ_BEW_RATE_CTRL    32'h00000102
`define DDRMC__REG_CMDQ_BEW_RATE_CTRL_SZ 22

`define DDRMC__REG_CMDQ_CTRL0    32'h00000103
`define DDRMC__REG_CMDQ_CTRL0_SZ 25

`define DDRMC__REG_CMDQ_CTRL1    32'h00000104
`define DDRMC__REG_CMDQ_CTRL1_SZ 25

`define DDRMC__REG_CMDQ_ISR_RATE_CTRL    32'h00000105
`define DDRMC__REG_CMDQ_ISR_RATE_CTRL_SZ 22

`define DDRMC__REG_CMDQ_ISW_RATE_CTRL    32'h00000106
`define DDRMC__REG_CMDQ_ISW_RATE_CTRL_SZ 22

`define DDRMC__REG_CMDQ_LLR_RATE_CTRL    32'h00000107
`define DDRMC__REG_CMDQ_LLR_RATE_CTRL_SZ 22

`define DDRMC__REG_COM_1    32'h00000108
`define DDRMC__REG_COM_1_SZ 27

`define DDRMC__REG_COM_2    32'h00000109
`define DDRMC__REG_COM_2_SZ 27

`define DDRMC__REG_COM_3    32'h0000010a
`define DDRMC__REG_COM_3_SZ 18

`define DDRMC__REG_CONFIG0    32'h0000010b
`define DDRMC__REG_CONFIG0_SZ 23

`define DDRMC__REG_CONFIG1    32'h0000010c
`define DDRMC__REG_CONFIG1_SZ 3

`define DDRMC__REG_CONFIG2    32'h0000010d
`define DDRMC__REG_CONFIG2_SZ 31

`define DDRMC__REG_CONFIG3    32'h0000010e
`define DDRMC__REG_CONFIG3_SZ 32

`define DDRMC__REG_CONFIG4    32'h0000010f
`define DDRMC__REG_CONFIG4_SZ 23

`define DDRMC__REG_DRAM_ARB    32'h00000110
`define DDRMC__REG_DRAM_ARB_SZ 13

`define DDRMC__REG_MRS_0    32'h00000111
`define DDRMC__REG_MRS_0_SZ 26

`define DDRMC__REG_MRS_1    32'h00000112
`define DDRMC__REG_MRS_1_SZ 32

`define DDRMC__REG_MRS_2    32'h00000113
`define DDRMC__REG_MRS_2_SZ 3

`define DDRMC__REG_MRS_7    32'h00000114
`define DDRMC__REG_MRS_7_SZ 8

`define DDRMC__REG_NSU0_PORT    32'h00000115
`define DDRMC__REG_NSU0_PORT_SZ 12

`define DDRMC__REG_NSU1_PORT    32'h00000116
`define DDRMC__REG_NSU1_PORT_SZ 12

`define DDRMC__REG_NSU2_PORT    32'h00000117
`define DDRMC__REG_NSU2_PORT_SZ 12

`define DDRMC__REG_NSU3_PORT    32'h00000118
`define DDRMC__REG_NSU3_PORT_SZ 12

`define DDRMC__REG_NSU_0_EGR    32'h00000119
`define DDRMC__REG_NSU_0_EGR_SZ 23

`define DDRMC__REG_NSU_0_ING    32'h0000011a
`define DDRMC__REG_NSU_0_ING_SZ 27

`define DDRMC__REG_NSU_0_R_EGR    32'h0000011b
`define DDRMC__REG_NSU_0_R_EGR_SZ 28

`define DDRMC__REG_NSU_0_W_EGR    32'h0000011c
`define DDRMC__REG_NSU_0_W_EGR_SZ 20

`define DDRMC__REG_NSU_1_EGR    32'h0000011d
`define DDRMC__REG_NSU_1_EGR_SZ 23

`define DDRMC__REG_NSU_1_ING    32'h0000011e
`define DDRMC__REG_NSU_1_ING_SZ 27

`define DDRMC__REG_NSU_1_R_EGR    32'h0000011f
`define DDRMC__REG_NSU_1_R_EGR_SZ 28

`define DDRMC__REG_NSU_1_W_EGR    32'h00000120
`define DDRMC__REG_NSU_1_W_EGR_SZ 20

`define DDRMC__REG_NSU_2_EGR    32'h00000121
`define DDRMC__REG_NSU_2_EGR_SZ 23

`define DDRMC__REG_NSU_2_ING    32'h00000122
`define DDRMC__REG_NSU_2_ING_SZ 27

`define DDRMC__REG_NSU_2_R_EGR    32'h00000123
`define DDRMC__REG_NSU_2_R_EGR_SZ 28

`define DDRMC__REG_NSU_2_W_EGR    32'h00000124
`define DDRMC__REG_NSU_2_W_EGR_SZ 20

`define DDRMC__REG_NSU_3_EGR    32'h00000125
`define DDRMC__REG_NSU_3_EGR_SZ 23

`define DDRMC__REG_NSU_3_ING    32'h00000126
`define DDRMC__REG_NSU_3_ING_SZ 27

`define DDRMC__REG_NSU_3_R_EGR    32'h00000127
`define DDRMC__REG_NSU_3_R_EGR_SZ 28

`define DDRMC__REG_NSU_3_W_EGR    32'h00000128
`define DDRMC__REG_NSU_3_W_EGR_SZ 20

`define DDRMC__REG_P0_BER_RATE_CTRL    32'h00000129
`define DDRMC__REG_P0_BER_RATE_CTRL_SZ 22

`define DDRMC__REG_P0_BEW_RATE_CTRL    32'h0000012a
`define DDRMC__REG_P0_BEW_RATE_CTRL_SZ 22

`define DDRMC__REG_P0_ISR_RATE_CTRL    32'h0000012b
`define DDRMC__REG_P0_ISR_RATE_CTRL_SZ 22

`define DDRMC__REG_P0_ISW_RATE_CTRL    32'h0000012c
`define DDRMC__REG_P0_ISW_RATE_CTRL_SZ 22

`define DDRMC__REG_P0_LLR_RATE_CTRL    32'h0000012d
`define DDRMC__REG_P0_LLR_RATE_CTRL_SZ 22

`define DDRMC__REG_P1_BER_RATE_CTRL    32'h0000012e
`define DDRMC__REG_P1_BER_RATE_CTRL_SZ 22

`define DDRMC__REG_P1_BEW_RATE_CTRL    32'h0000012f
`define DDRMC__REG_P1_BEW_RATE_CTRL_SZ 22

`define DDRMC__REG_P1_ISR_RATE_CTRL    32'h00000130
`define DDRMC__REG_P1_ISR_RATE_CTRL_SZ 22

`define DDRMC__REG_P1_ISW_RATE_CTRL    32'h00000131
`define DDRMC__REG_P1_ISW_RATE_CTRL_SZ 22

`define DDRMC__REG_P1_LLR_RATE_CTRL    32'h00000132
`define DDRMC__REG_P1_LLR_RATE_CTRL_SZ 22

`define DDRMC__REG_P2_BER_RATE_CTRL    32'h00000133
`define DDRMC__REG_P2_BER_RATE_CTRL_SZ 22

`define DDRMC__REG_P2_BEW_RATE_CTRL    32'h00000134
`define DDRMC__REG_P2_BEW_RATE_CTRL_SZ 22

`define DDRMC__REG_P2_ISR_RATE_CTRL    32'h00000135
`define DDRMC__REG_P2_ISR_RATE_CTRL_SZ 22

`define DDRMC__REG_P2_ISW_RATE_CTRL    32'h00000136
`define DDRMC__REG_P2_ISW_RATE_CTRL_SZ 22

`define DDRMC__REG_P2_LLR_RATE_CTRL    32'h00000137
`define DDRMC__REG_P2_LLR_RATE_CTRL_SZ 22

`define DDRMC__REG_P3_BER_RATE_CTRL    32'h00000138
`define DDRMC__REG_P3_BER_RATE_CTRL_SZ 22

`define DDRMC__REG_P3_BEW_RATE_CTRL    32'h00000139
`define DDRMC__REG_P3_BEW_RATE_CTRL_SZ 22

`define DDRMC__REG_P3_ISR_RATE_CTRL    32'h0000013a
`define DDRMC__REG_P3_ISR_RATE_CTRL_SZ 22

`define DDRMC__REG_P3_ISW_RATE_CTRL    32'h0000013b
`define DDRMC__REG_P3_ISW_RATE_CTRL_SZ 22

`define DDRMC__REG_P3_LLR_RATE_CTRL    32'h0000013c
`define DDRMC__REG_P3_LLR_RATE_CTRL_SZ 22

`define DDRMC__REG_PINOUT    32'h0000013d
`define DDRMC__REG_PINOUT_SZ 10

`define DDRMC__REG_PT_CONFIG    32'h0000013e
`define DDRMC__REG_PT_CONFIG_SZ 20

`define DDRMC__REG_QOS0    32'h0000013f
`define DDRMC__REG_QOS0_SZ 28

`define DDRMC__REG_QOS1    32'h00000140
`define DDRMC__REG_QOS1_SZ 30

`define DDRMC__REG_QOS2    32'h00000141
`define DDRMC__REG_QOS2_SZ 20

`define DDRMC__REG_QOS_RATE_CTRL_SCALE    32'h00000142
`define DDRMC__REG_QOS_RATE_CTRL_SCALE_SZ 25

`define DDRMC__REG_QOS_TIMEOUT0    32'h00000143
`define DDRMC__REG_QOS_TIMEOUT0_SZ 25

`define DDRMC__REG_QOS_TIMEOUT1    32'h00000144
`define DDRMC__REG_QOS_TIMEOUT1_SZ 32

`define DDRMC__REG_QOS_TIMEOUT2    32'h00000145
`define DDRMC__REG_QOS_TIMEOUT2_SZ 8

`define DDRMC__REG_RATE_CTRL_SCALE    32'h00000146
`define DDRMC__REG_RATE_CTRL_SCALE_SZ 25

`define DDRMC__REG_RD_CONFIG    32'h00000147
`define DDRMC__REG_RD_CONFIG_SZ 30

`define DDRMC__REG_RD_DRR_TKN_P0    32'h00000148
`define DDRMC__REG_RD_DRR_TKN_P0_SZ 24

`define DDRMC__REG_RD_DRR_TKN_P1    32'h00000149
`define DDRMC__REG_RD_DRR_TKN_P1_SZ 24

`define DDRMC__REG_RD_DRR_TKN_P2    32'h0000014a
`define DDRMC__REG_RD_DRR_TKN_P2_SZ 24

`define DDRMC__REG_RD_DRR_TKN_P3    32'h0000014b
`define DDRMC__REG_RD_DRR_TKN_P3_SZ 24

`define DDRMC__REG_REF_0    32'h0000014c
`define DDRMC__REG_REF_0_SZ 2

`define DDRMC__REG_REF_1    32'h0000014d
`define DDRMC__REG_REF_1_SZ 32

`define DDRMC__REG_REF_2    32'h0000014e
`define DDRMC__REG_REF_2_SZ 2

`define DDRMC__REG_REF_3    32'h0000014f
`define DDRMC__REG_REF_3_SZ 16

`define DDRMC__REG_RETRY_0    32'h00000150
`define DDRMC__REG_RETRY_0_SZ 29

`define DDRMC__REG_RETRY_1    32'h00000151
`define DDRMC__REG_RETRY_1_SZ 30

`define DDRMC__REG_SAFE_CONFIG0    32'h00000152
`define DDRMC__REG_SAFE_CONFIG0_SZ 32

`define DDRMC__REG_SAFE_CONFIG1    32'h00000153
`define DDRMC__REG_SAFE_CONFIG1_SZ 32

`define DDRMC__REG_SAFE_CONFIG2    32'h00000154
`define DDRMC__REG_SAFE_CONFIG2_SZ 32

`define DDRMC__REG_SAFE_CONFIG3    32'h00000155
`define DDRMC__REG_SAFE_CONFIG3_SZ 28

`define DDRMC__REG_SAFE_CONFIG4    32'h00000156
`define DDRMC__REG_SAFE_CONFIG4_SZ 31

`define DDRMC__REG_SAFE_CONFIG5    32'h00000157
`define DDRMC__REG_SAFE_CONFIG5_SZ 32

`define DDRMC__REG_SAFE_CONFIG6    32'h00000158
`define DDRMC__REG_SAFE_CONFIG6_SZ 26

`define DDRMC__REG_SAFE_CONFIG7    32'h00000159
`define DDRMC__REG_SAFE_CONFIG7_SZ 30

`define DDRMC__REG_SAFE_CONFIG8    32'h0000015a
`define DDRMC__REG_SAFE_CONFIG8_SZ 32

`define DDRMC__REG_SCRUB0    32'h0000015b
`define DDRMC__REG_SCRUB0_SZ 32

`define DDRMC__REG_SCRUB1    32'h0000015c
`define DDRMC__REG_SCRUB1_SZ 32

`define DDRMC__REG_SCRUB8    32'h0000015d
`define DDRMC__REG_SCRUB8_SZ 2

`define DDRMC__REG_SCRUB9    32'h0000015e
`define DDRMC__REG_SCRUB9_SZ 1

`define DDRMC__REG_TXN_CONFIG    32'h0000015f
`define DDRMC__REG_TXN_CONFIG_SZ 20

`define DDRMC__REG_WR_CONFIG    32'h00000160
`define DDRMC__REG_WR_CONFIG_SZ 32

`define DDRMC__REG_WR_DRR_TKN_P0    32'h00000161
`define DDRMC__REG_WR_DRR_TKN_P0_SZ 16

`define DDRMC__REG_WR_DRR_TKN_P1    32'h00000162
`define DDRMC__REG_WR_DRR_TKN_P1_SZ 16

`define DDRMC__REG_WR_DRR_TKN_P2    32'h00000163
`define DDRMC__REG_WR_DRR_TKN_P2_SZ 16

`define DDRMC__REG_WR_DRR_TKN_P3    32'h00000164
`define DDRMC__REG_WR_DRR_TKN_P3_SZ 16

`define DDRMC__SEQ_ADDR_DEFAULT    32'h00000165
`define DDRMC__SEQ_ADDR_DEFAULT_SZ 1

`define DDRMC__SEQ_BA_DEFAULT    32'h00000166
`define DDRMC__SEQ_BA_DEFAULT_SZ 1

`define DDRMC__SEQ_BG_DEFAULT    32'h00000167
`define DDRMC__SEQ_BG_DEFAULT_SZ 1

`define DDRMC__SEQ_CBIT_DEFAULT    32'h00000168
`define DDRMC__SEQ_CBIT_DEFAULT_SZ 1

`define DDRMC__SEQ_CK_CAL    32'h00000169
`define DDRMC__SEQ_CK_CAL_SZ 16

`define DDRMC__SEQ_CMD_DEFAULT    32'h0000016a
`define DDRMC__SEQ_CMD_DEFAULT_SZ 7

`define DDRMC__SEQ_CMD_POR    32'h0000016b
`define DDRMC__SEQ_CMD_POR_SZ 7

`define DDRMC__SEQ_DQS_DEFAULT    32'h0000016c
`define DDRMC__SEQ_DQS_DEFAULT_SZ 3

`define DDRMC__SEQ_DQ_DEFAULT    32'h0000016d
`define DDRMC__SEQ_DQ_DEFAULT_SZ 5

`define DDRMC__SEQ_INIT_ADDR0    32'h0000016e
`define DDRMC__SEQ_INIT_ADDR0_SZ 28

`define DDRMC__SEQ_INIT_ADDR1    32'h0000016f
`define DDRMC__SEQ_INIT_ADDR1_SZ 28

`define DDRMC__SEQ_INIT_ADDR10    32'h00000170
`define DDRMC__SEQ_INIT_ADDR10_SZ 28

`define DDRMC__SEQ_INIT_ADDR11    32'h00000171
`define DDRMC__SEQ_INIT_ADDR11_SZ 28

`define DDRMC__SEQ_INIT_ADDR12    32'h00000172
`define DDRMC__SEQ_INIT_ADDR12_SZ 28

`define DDRMC__SEQ_INIT_ADDR13    32'h00000173
`define DDRMC__SEQ_INIT_ADDR13_SZ 28

`define DDRMC__SEQ_INIT_ADDR14    32'h00000174
`define DDRMC__SEQ_INIT_ADDR14_SZ 28

`define DDRMC__SEQ_INIT_ADDR15    32'h00000175
`define DDRMC__SEQ_INIT_ADDR15_SZ 28

`define DDRMC__SEQ_INIT_ADDR16    32'h00000176
`define DDRMC__SEQ_INIT_ADDR16_SZ 28

`define DDRMC__SEQ_INIT_ADDR17    32'h00000177
`define DDRMC__SEQ_INIT_ADDR17_SZ 28

`define DDRMC__SEQ_INIT_ADDR18    32'h00000178
`define DDRMC__SEQ_INIT_ADDR18_SZ 28

`define DDRMC__SEQ_INIT_ADDR19    32'h00000179
`define DDRMC__SEQ_INIT_ADDR19_SZ 28

`define DDRMC__SEQ_INIT_ADDR2    32'h0000017a
`define DDRMC__SEQ_INIT_ADDR2_SZ 28

`define DDRMC__SEQ_INIT_ADDR20    32'h0000017b
`define DDRMC__SEQ_INIT_ADDR20_SZ 28

`define DDRMC__SEQ_INIT_ADDR21    32'h0000017c
`define DDRMC__SEQ_INIT_ADDR21_SZ 28

`define DDRMC__SEQ_INIT_ADDR22    32'h0000017d
`define DDRMC__SEQ_INIT_ADDR22_SZ 28

`define DDRMC__SEQ_INIT_ADDR23    32'h0000017e
`define DDRMC__SEQ_INIT_ADDR23_SZ 28

`define DDRMC__SEQ_INIT_ADDR24    32'h0000017f
`define DDRMC__SEQ_INIT_ADDR24_SZ 28

`define DDRMC__SEQ_INIT_ADDR25    32'h00000180
`define DDRMC__SEQ_INIT_ADDR25_SZ 28

`define DDRMC__SEQ_INIT_ADDR26    32'h00000181
`define DDRMC__SEQ_INIT_ADDR26_SZ 28

`define DDRMC__SEQ_INIT_ADDR27    32'h00000182
`define DDRMC__SEQ_INIT_ADDR27_SZ 28

`define DDRMC__SEQ_INIT_ADDR28    32'h00000183
`define DDRMC__SEQ_INIT_ADDR28_SZ 28

`define DDRMC__SEQ_INIT_ADDR29    32'h00000184
`define DDRMC__SEQ_INIT_ADDR29_SZ 28

`define DDRMC__SEQ_INIT_ADDR3    32'h00000185
`define DDRMC__SEQ_INIT_ADDR3_SZ 28

`define DDRMC__SEQ_INIT_ADDR30    32'h00000186
`define DDRMC__SEQ_INIT_ADDR30_SZ 28

`define DDRMC__SEQ_INIT_ADDR31    32'h00000187
`define DDRMC__SEQ_INIT_ADDR31_SZ 28

`define DDRMC__SEQ_INIT_ADDR32    32'h00000188
`define DDRMC__SEQ_INIT_ADDR32_SZ 28

`define DDRMC__SEQ_INIT_ADDR33    32'h00000189
`define DDRMC__SEQ_INIT_ADDR33_SZ 28

`define DDRMC__SEQ_INIT_ADDR34    32'h0000018a
`define DDRMC__SEQ_INIT_ADDR34_SZ 28

`define DDRMC__SEQ_INIT_ADDR35    32'h0000018b
`define DDRMC__SEQ_INIT_ADDR35_SZ 28

`define DDRMC__SEQ_INIT_ADDR36    32'h0000018c
`define DDRMC__SEQ_INIT_ADDR36_SZ 28

`define DDRMC__SEQ_INIT_ADDR37    32'h0000018d
`define DDRMC__SEQ_INIT_ADDR37_SZ 28

`define DDRMC__SEQ_INIT_ADDR38    32'h0000018e
`define DDRMC__SEQ_INIT_ADDR38_SZ 28

`define DDRMC__SEQ_INIT_ADDR39    32'h0000018f
`define DDRMC__SEQ_INIT_ADDR39_SZ 28

`define DDRMC__SEQ_INIT_ADDR4    32'h00000190
`define DDRMC__SEQ_INIT_ADDR4_SZ 28

`define DDRMC__SEQ_INIT_ADDR40    32'h00000191
`define DDRMC__SEQ_INIT_ADDR40_SZ 28

`define DDRMC__SEQ_INIT_ADDR41    32'h00000192
`define DDRMC__SEQ_INIT_ADDR41_SZ 28

`define DDRMC__SEQ_INIT_ADDR42    32'h00000193
`define DDRMC__SEQ_INIT_ADDR42_SZ 28

`define DDRMC__SEQ_INIT_ADDR43    32'h00000194
`define DDRMC__SEQ_INIT_ADDR43_SZ 28

`define DDRMC__SEQ_INIT_ADDR44    32'h00000195
`define DDRMC__SEQ_INIT_ADDR44_SZ 28

`define DDRMC__SEQ_INIT_ADDR45    32'h00000196
`define DDRMC__SEQ_INIT_ADDR45_SZ 28

`define DDRMC__SEQ_INIT_ADDR46    32'h00000197
`define DDRMC__SEQ_INIT_ADDR46_SZ 28

`define DDRMC__SEQ_INIT_ADDR47    32'h00000198
`define DDRMC__SEQ_INIT_ADDR47_SZ 28

`define DDRMC__SEQ_INIT_ADDR48    32'h00000199
`define DDRMC__SEQ_INIT_ADDR48_SZ 28

`define DDRMC__SEQ_INIT_ADDR49    32'h0000019a
`define DDRMC__SEQ_INIT_ADDR49_SZ 28

`define DDRMC__SEQ_INIT_ADDR5    32'h0000019b
`define DDRMC__SEQ_INIT_ADDR5_SZ 28

`define DDRMC__SEQ_INIT_ADDR50    32'h0000019c
`define DDRMC__SEQ_INIT_ADDR50_SZ 28

`define DDRMC__SEQ_INIT_ADDR51    32'h0000019d
`define DDRMC__SEQ_INIT_ADDR51_SZ 28

`define DDRMC__SEQ_INIT_ADDR52    32'h0000019e
`define DDRMC__SEQ_INIT_ADDR52_SZ 28

`define DDRMC__SEQ_INIT_ADDR53    32'h0000019f
`define DDRMC__SEQ_INIT_ADDR53_SZ 28

`define DDRMC__SEQ_INIT_ADDR54    32'h000001a0
`define DDRMC__SEQ_INIT_ADDR54_SZ 28

`define DDRMC__SEQ_INIT_ADDR55    32'h000001a1
`define DDRMC__SEQ_INIT_ADDR55_SZ 28

`define DDRMC__SEQ_INIT_ADDR56    32'h000001a2
`define DDRMC__SEQ_INIT_ADDR56_SZ 28

`define DDRMC__SEQ_INIT_ADDR57    32'h000001a3
`define DDRMC__SEQ_INIT_ADDR57_SZ 28

`define DDRMC__SEQ_INIT_ADDR58    32'h000001a4
`define DDRMC__SEQ_INIT_ADDR58_SZ 28

`define DDRMC__SEQ_INIT_ADDR59    32'h000001a5
`define DDRMC__SEQ_INIT_ADDR59_SZ 28

`define DDRMC__SEQ_INIT_ADDR6    32'h000001a6
`define DDRMC__SEQ_INIT_ADDR6_SZ 28

`define DDRMC__SEQ_INIT_ADDR60    32'h000001a7
`define DDRMC__SEQ_INIT_ADDR60_SZ 28

`define DDRMC__SEQ_INIT_ADDR61    32'h000001a8
`define DDRMC__SEQ_INIT_ADDR61_SZ 28

`define DDRMC__SEQ_INIT_ADDR62    32'h000001a9
`define DDRMC__SEQ_INIT_ADDR62_SZ 28

`define DDRMC__SEQ_INIT_ADDR63    32'h000001aa
`define DDRMC__SEQ_INIT_ADDR63_SZ 28

`define DDRMC__SEQ_INIT_ADDR64    32'h000001ab
`define DDRMC__SEQ_INIT_ADDR64_SZ 28

`define DDRMC__SEQ_INIT_ADDR65    32'h000001ac
`define DDRMC__SEQ_INIT_ADDR65_SZ 28

`define DDRMC__SEQ_INIT_ADDR66    32'h000001ad
`define DDRMC__SEQ_INIT_ADDR66_SZ 28

`define DDRMC__SEQ_INIT_ADDR67    32'h000001ae
`define DDRMC__SEQ_INIT_ADDR67_SZ 28

`define DDRMC__SEQ_INIT_ADDR68    32'h000001af
`define DDRMC__SEQ_INIT_ADDR68_SZ 28

`define DDRMC__SEQ_INIT_ADDR69    32'h000001b0
`define DDRMC__SEQ_INIT_ADDR69_SZ 28

`define DDRMC__SEQ_INIT_ADDR7    32'h000001b1
`define DDRMC__SEQ_INIT_ADDR7_SZ 28

`define DDRMC__SEQ_INIT_ADDR70    32'h000001b2
`define DDRMC__SEQ_INIT_ADDR70_SZ 28

`define DDRMC__SEQ_INIT_ADDR71    32'h000001b3
`define DDRMC__SEQ_INIT_ADDR71_SZ 28

`define DDRMC__SEQ_INIT_ADDR72    32'h000001b4
`define DDRMC__SEQ_INIT_ADDR72_SZ 28

`define DDRMC__SEQ_INIT_ADDR73    32'h000001b5
`define DDRMC__SEQ_INIT_ADDR73_SZ 28

`define DDRMC__SEQ_INIT_ADDR74    32'h000001b6
`define DDRMC__SEQ_INIT_ADDR74_SZ 28

`define DDRMC__SEQ_INIT_ADDR75    32'h000001b7
`define DDRMC__SEQ_INIT_ADDR75_SZ 28

`define DDRMC__SEQ_INIT_ADDR76    32'h000001b8
`define DDRMC__SEQ_INIT_ADDR76_SZ 28

`define DDRMC__SEQ_INIT_ADDR77    32'h000001b9
`define DDRMC__SEQ_INIT_ADDR77_SZ 28

`define DDRMC__SEQ_INIT_ADDR78    32'h000001ba
`define DDRMC__SEQ_INIT_ADDR78_SZ 28

`define DDRMC__SEQ_INIT_ADDR79    32'h000001bb
`define DDRMC__SEQ_INIT_ADDR79_SZ 28

`define DDRMC__SEQ_INIT_ADDR8    32'h000001bc
`define DDRMC__SEQ_INIT_ADDR8_SZ 28

`define DDRMC__SEQ_INIT_ADDR80    32'h000001bd
`define DDRMC__SEQ_INIT_ADDR80_SZ 28

`define DDRMC__SEQ_INIT_ADDR81    32'h000001be
`define DDRMC__SEQ_INIT_ADDR81_SZ 28

`define DDRMC__SEQ_INIT_ADDR82    32'h000001bf
`define DDRMC__SEQ_INIT_ADDR82_SZ 28

`define DDRMC__SEQ_INIT_ADDR83    32'h000001c0
`define DDRMC__SEQ_INIT_ADDR83_SZ 28

`define DDRMC__SEQ_INIT_ADDR84    32'h000001c1
`define DDRMC__SEQ_INIT_ADDR84_SZ 28

`define DDRMC__SEQ_INIT_ADDR85    32'h000001c2
`define DDRMC__SEQ_INIT_ADDR85_SZ 28

`define DDRMC__SEQ_INIT_ADDR86    32'h000001c3
`define DDRMC__SEQ_INIT_ADDR86_SZ 28

`define DDRMC__SEQ_INIT_ADDR87    32'h000001c4
`define DDRMC__SEQ_INIT_ADDR87_SZ 28

`define DDRMC__SEQ_INIT_ADDR88    32'h000001c5
`define DDRMC__SEQ_INIT_ADDR88_SZ 28

`define DDRMC__SEQ_INIT_ADDR89    32'h000001c6
`define DDRMC__SEQ_INIT_ADDR89_SZ 28

`define DDRMC__SEQ_INIT_ADDR9    32'h000001c7
`define DDRMC__SEQ_INIT_ADDR9_SZ 28

`define DDRMC__SEQ_INIT_ADDR90    32'h000001c8
`define DDRMC__SEQ_INIT_ADDR90_SZ 28

`define DDRMC__SEQ_INIT_ADDR91    32'h000001c9
`define DDRMC__SEQ_INIT_ADDR91_SZ 28

`define DDRMC__SEQ_INIT_ADDR92    32'h000001ca
`define DDRMC__SEQ_INIT_ADDR92_SZ 28

`define DDRMC__SEQ_INIT_ADDR93    32'h000001cb
`define DDRMC__SEQ_INIT_ADDR93_SZ 28

`define DDRMC__SEQ_INIT_ADDR94    32'h000001cc
`define DDRMC__SEQ_INIT_ADDR94_SZ 28

`define DDRMC__SEQ_INIT_ADDR95    32'h000001cd
`define DDRMC__SEQ_INIT_ADDR95_SZ 28

`define DDRMC__SEQ_INIT_ADDR96    32'h000001ce
`define DDRMC__SEQ_INIT_ADDR96_SZ 28

`define DDRMC__SEQ_INIT_ADDR97    32'h000001cf
`define DDRMC__SEQ_INIT_ADDR97_SZ 28

`define DDRMC__SEQ_INIT_ADDR98    32'h000001d0
`define DDRMC__SEQ_INIT_ADDR98_SZ 28

`define DDRMC__SEQ_INIT_ADDR99    32'h000001d1
`define DDRMC__SEQ_INIT_ADDR99_SZ 28

`define DDRMC__SEQ_INIT_CMD0    32'h000001d2
`define DDRMC__SEQ_INIT_CMD0_SZ 32

`define DDRMC__SEQ_INIT_CMD1    32'h000001d3
`define DDRMC__SEQ_INIT_CMD1_SZ 32

`define DDRMC__SEQ_INIT_CMD10    32'h000001d4
`define DDRMC__SEQ_INIT_CMD10_SZ 32

`define DDRMC__SEQ_INIT_CMD11    32'h000001d5
`define DDRMC__SEQ_INIT_CMD11_SZ 32

`define DDRMC__SEQ_INIT_CMD12    32'h000001d6
`define DDRMC__SEQ_INIT_CMD12_SZ 32

`define DDRMC__SEQ_INIT_CMD13    32'h000001d7
`define DDRMC__SEQ_INIT_CMD13_SZ 32

`define DDRMC__SEQ_INIT_CMD14    32'h000001d8
`define DDRMC__SEQ_INIT_CMD14_SZ 32

`define DDRMC__SEQ_INIT_CMD15    32'h000001d9
`define DDRMC__SEQ_INIT_CMD15_SZ 32

`define DDRMC__SEQ_INIT_CMD16    32'h000001da
`define DDRMC__SEQ_INIT_CMD16_SZ 32

`define DDRMC__SEQ_INIT_CMD17    32'h000001db
`define DDRMC__SEQ_INIT_CMD17_SZ 32

`define DDRMC__SEQ_INIT_CMD18    32'h000001dc
`define DDRMC__SEQ_INIT_CMD18_SZ 32

`define DDRMC__SEQ_INIT_CMD19    32'h000001dd
`define DDRMC__SEQ_INIT_CMD19_SZ 32

`define DDRMC__SEQ_INIT_CMD2    32'h000001de
`define DDRMC__SEQ_INIT_CMD2_SZ 32

`define DDRMC__SEQ_INIT_CMD20    32'h000001df
`define DDRMC__SEQ_INIT_CMD20_SZ 32

`define DDRMC__SEQ_INIT_CMD21    32'h000001e0
`define DDRMC__SEQ_INIT_CMD21_SZ 32

`define DDRMC__SEQ_INIT_CMD22    32'h000001e1
`define DDRMC__SEQ_INIT_CMD22_SZ 32

`define DDRMC__SEQ_INIT_CMD23    32'h000001e2
`define DDRMC__SEQ_INIT_CMD23_SZ 32

`define DDRMC__SEQ_INIT_CMD24    32'h000001e3
`define DDRMC__SEQ_INIT_CMD24_SZ 32

`define DDRMC__SEQ_INIT_CMD25    32'h000001e4
`define DDRMC__SEQ_INIT_CMD25_SZ 32

`define DDRMC__SEQ_INIT_CMD26    32'h000001e5
`define DDRMC__SEQ_INIT_CMD26_SZ 32

`define DDRMC__SEQ_INIT_CMD27    32'h000001e6
`define DDRMC__SEQ_INIT_CMD27_SZ 32

`define DDRMC__SEQ_INIT_CMD28    32'h000001e7
`define DDRMC__SEQ_INIT_CMD28_SZ 32

`define DDRMC__SEQ_INIT_CMD29    32'h000001e8
`define DDRMC__SEQ_INIT_CMD29_SZ 32

`define DDRMC__SEQ_INIT_CMD3    32'h000001e9
`define DDRMC__SEQ_INIT_CMD3_SZ 32

`define DDRMC__SEQ_INIT_CMD30    32'h000001ea
`define DDRMC__SEQ_INIT_CMD30_SZ 32

`define DDRMC__SEQ_INIT_CMD31    32'h000001eb
`define DDRMC__SEQ_INIT_CMD31_SZ 32

`define DDRMC__SEQ_INIT_CMD32    32'h000001ec
`define DDRMC__SEQ_INIT_CMD32_SZ 32

`define DDRMC__SEQ_INIT_CMD33    32'h000001ed
`define DDRMC__SEQ_INIT_CMD33_SZ 32

`define DDRMC__SEQ_INIT_CMD34    32'h000001ee
`define DDRMC__SEQ_INIT_CMD34_SZ 32

`define DDRMC__SEQ_INIT_CMD35    32'h000001ef
`define DDRMC__SEQ_INIT_CMD35_SZ 32

`define DDRMC__SEQ_INIT_CMD36    32'h000001f0
`define DDRMC__SEQ_INIT_CMD36_SZ 32

`define DDRMC__SEQ_INIT_CMD37    32'h000001f1
`define DDRMC__SEQ_INIT_CMD37_SZ 32

`define DDRMC__SEQ_INIT_CMD38    32'h000001f2
`define DDRMC__SEQ_INIT_CMD38_SZ 32

`define DDRMC__SEQ_INIT_CMD39    32'h000001f3
`define DDRMC__SEQ_INIT_CMD39_SZ 32

`define DDRMC__SEQ_INIT_CMD4    32'h000001f4
`define DDRMC__SEQ_INIT_CMD4_SZ 32

`define DDRMC__SEQ_INIT_CMD40    32'h000001f5
`define DDRMC__SEQ_INIT_CMD40_SZ 32

`define DDRMC__SEQ_INIT_CMD41    32'h000001f6
`define DDRMC__SEQ_INIT_CMD41_SZ 32

`define DDRMC__SEQ_INIT_CMD42    32'h000001f7
`define DDRMC__SEQ_INIT_CMD42_SZ 32

`define DDRMC__SEQ_INIT_CMD43    32'h000001f8
`define DDRMC__SEQ_INIT_CMD43_SZ 32

`define DDRMC__SEQ_INIT_CMD44    32'h000001f9
`define DDRMC__SEQ_INIT_CMD44_SZ 32

`define DDRMC__SEQ_INIT_CMD45    32'h000001fa
`define DDRMC__SEQ_INIT_CMD45_SZ 32

`define DDRMC__SEQ_INIT_CMD46    32'h000001fb
`define DDRMC__SEQ_INIT_CMD46_SZ 32

`define DDRMC__SEQ_INIT_CMD47    32'h000001fc
`define DDRMC__SEQ_INIT_CMD47_SZ 32

`define DDRMC__SEQ_INIT_CMD48    32'h000001fd
`define DDRMC__SEQ_INIT_CMD48_SZ 32

`define DDRMC__SEQ_INIT_CMD49    32'h000001fe
`define DDRMC__SEQ_INIT_CMD49_SZ 32

`define DDRMC__SEQ_INIT_CMD5    32'h000001ff
`define DDRMC__SEQ_INIT_CMD5_SZ 32

`define DDRMC__SEQ_INIT_CMD50    32'h00000200
`define DDRMC__SEQ_INIT_CMD50_SZ 32

`define DDRMC__SEQ_INIT_CMD51    32'h00000201
`define DDRMC__SEQ_INIT_CMD51_SZ 32

`define DDRMC__SEQ_INIT_CMD52    32'h00000202
`define DDRMC__SEQ_INIT_CMD52_SZ 32

`define DDRMC__SEQ_INIT_CMD53    32'h00000203
`define DDRMC__SEQ_INIT_CMD53_SZ 32

`define DDRMC__SEQ_INIT_CMD54    32'h00000204
`define DDRMC__SEQ_INIT_CMD54_SZ 32

`define DDRMC__SEQ_INIT_CMD55    32'h00000205
`define DDRMC__SEQ_INIT_CMD55_SZ 32

`define DDRMC__SEQ_INIT_CMD56    32'h00000206
`define DDRMC__SEQ_INIT_CMD56_SZ 32

`define DDRMC__SEQ_INIT_CMD57    32'h00000207
`define DDRMC__SEQ_INIT_CMD57_SZ 32

`define DDRMC__SEQ_INIT_CMD58    32'h00000208
`define DDRMC__SEQ_INIT_CMD58_SZ 32

`define DDRMC__SEQ_INIT_CMD59    32'h00000209
`define DDRMC__SEQ_INIT_CMD59_SZ 32

`define DDRMC__SEQ_INIT_CMD6    32'h0000020a
`define DDRMC__SEQ_INIT_CMD6_SZ 32

`define DDRMC__SEQ_INIT_CMD60    32'h0000020b
`define DDRMC__SEQ_INIT_CMD60_SZ 32

`define DDRMC__SEQ_INIT_CMD61    32'h0000020c
`define DDRMC__SEQ_INIT_CMD61_SZ 32

`define DDRMC__SEQ_INIT_CMD62    32'h0000020d
`define DDRMC__SEQ_INIT_CMD62_SZ 32

`define DDRMC__SEQ_INIT_CMD63    32'h0000020e
`define DDRMC__SEQ_INIT_CMD63_SZ 32

`define DDRMC__SEQ_INIT_CMD64    32'h0000020f
`define DDRMC__SEQ_INIT_CMD64_SZ 32

`define DDRMC__SEQ_INIT_CMD65    32'h00000210
`define DDRMC__SEQ_INIT_CMD65_SZ 32

`define DDRMC__SEQ_INIT_CMD66    32'h00000211
`define DDRMC__SEQ_INIT_CMD66_SZ 32

`define DDRMC__SEQ_INIT_CMD67    32'h00000212
`define DDRMC__SEQ_INIT_CMD67_SZ 32

`define DDRMC__SEQ_INIT_CMD68    32'h00000213
`define DDRMC__SEQ_INIT_CMD68_SZ 32

`define DDRMC__SEQ_INIT_CMD69    32'h00000214
`define DDRMC__SEQ_INIT_CMD69_SZ 32

`define DDRMC__SEQ_INIT_CMD7    32'h00000215
`define DDRMC__SEQ_INIT_CMD7_SZ 32

`define DDRMC__SEQ_INIT_CMD70    32'h00000216
`define DDRMC__SEQ_INIT_CMD70_SZ 32

`define DDRMC__SEQ_INIT_CMD71    32'h00000217
`define DDRMC__SEQ_INIT_CMD71_SZ 32

`define DDRMC__SEQ_INIT_CMD72    32'h00000218
`define DDRMC__SEQ_INIT_CMD72_SZ 32

`define DDRMC__SEQ_INIT_CMD73    32'h00000219
`define DDRMC__SEQ_INIT_CMD73_SZ 32

`define DDRMC__SEQ_INIT_CMD74    32'h0000021a
`define DDRMC__SEQ_INIT_CMD74_SZ 32

`define DDRMC__SEQ_INIT_CMD75    32'h0000021b
`define DDRMC__SEQ_INIT_CMD75_SZ 32

`define DDRMC__SEQ_INIT_CMD76    32'h0000021c
`define DDRMC__SEQ_INIT_CMD76_SZ 32

`define DDRMC__SEQ_INIT_CMD77    32'h0000021d
`define DDRMC__SEQ_INIT_CMD77_SZ 32

`define DDRMC__SEQ_INIT_CMD78    32'h0000021e
`define DDRMC__SEQ_INIT_CMD78_SZ 32

`define DDRMC__SEQ_INIT_CMD79    32'h0000021f
`define DDRMC__SEQ_INIT_CMD79_SZ 32

`define DDRMC__SEQ_INIT_CMD8    32'h00000220
`define DDRMC__SEQ_INIT_CMD8_SZ 32

`define DDRMC__SEQ_INIT_CMD80    32'h00000221
`define DDRMC__SEQ_INIT_CMD80_SZ 32

`define DDRMC__SEQ_INIT_CMD81    32'h00000222
`define DDRMC__SEQ_INIT_CMD81_SZ 32

`define DDRMC__SEQ_INIT_CMD82    32'h00000223
`define DDRMC__SEQ_INIT_CMD82_SZ 32

`define DDRMC__SEQ_INIT_CMD83    32'h00000224
`define DDRMC__SEQ_INIT_CMD83_SZ 32

`define DDRMC__SEQ_INIT_CMD84    32'h00000225
`define DDRMC__SEQ_INIT_CMD84_SZ 32

`define DDRMC__SEQ_INIT_CMD85    32'h00000226
`define DDRMC__SEQ_INIT_CMD85_SZ 32

`define DDRMC__SEQ_INIT_CMD86    32'h00000227
`define DDRMC__SEQ_INIT_CMD86_SZ 32

`define DDRMC__SEQ_INIT_CMD87    32'h00000228
`define DDRMC__SEQ_INIT_CMD87_SZ 32

`define DDRMC__SEQ_INIT_CMD88    32'h00000229
`define DDRMC__SEQ_INIT_CMD88_SZ 32

`define DDRMC__SEQ_INIT_CMD89    32'h0000022a
`define DDRMC__SEQ_INIT_CMD89_SZ 32

`define DDRMC__SEQ_INIT_CMD9    32'h0000022b
`define DDRMC__SEQ_INIT_CMD9_SZ 32

`define DDRMC__SEQ_INIT_CMD90    32'h0000022c
`define DDRMC__SEQ_INIT_CMD90_SZ 32

`define DDRMC__SEQ_INIT_CMD91    32'h0000022d
`define DDRMC__SEQ_INIT_CMD91_SZ 32

`define DDRMC__SEQ_INIT_CMD92    32'h0000022e
`define DDRMC__SEQ_INIT_CMD92_SZ 32

`define DDRMC__SEQ_INIT_CMD93    32'h0000022f
`define DDRMC__SEQ_INIT_CMD93_SZ 32

`define DDRMC__SEQ_INIT_CMD94    32'h00000230
`define DDRMC__SEQ_INIT_CMD94_SZ 32

`define DDRMC__SEQ_INIT_CMD95    32'h00000231
`define DDRMC__SEQ_INIT_CMD95_SZ 32

`define DDRMC__SEQ_INIT_CMD96    32'h00000232
`define DDRMC__SEQ_INIT_CMD96_SZ 32

`define DDRMC__SEQ_INIT_CMD97    32'h00000233
`define DDRMC__SEQ_INIT_CMD97_SZ 32

`define DDRMC__SEQ_INIT_CMD98    32'h00000234
`define DDRMC__SEQ_INIT_CMD98_SZ 32

`define DDRMC__SEQ_INIT_CMD99    32'h00000235
`define DDRMC__SEQ_INIT_CMD99_SZ 32

`define DDRMC__SEQ_INIT_CMD_SET    32'h00000236
`define DDRMC__SEQ_INIT_CMD_SET_SZ 9

`define DDRMC__SEQ_INIT_CMD_VALID    32'h00000237
`define DDRMC__SEQ_INIT_CMD_VALID_SZ 7

`define DDRMC__SEQ_INIT_CNTRL0    32'h00000238
`define DDRMC__SEQ_INIT_CNTRL0_SZ 10

`define DDRMC__SEQ_INIT_CNTRL1    32'h00000239
`define DDRMC__SEQ_INIT_CNTRL1_SZ 10

`define DDRMC__SEQ_INIT_CNTRL10    32'h0000023a
`define DDRMC__SEQ_INIT_CNTRL10_SZ 10

`define DDRMC__SEQ_INIT_CNTRL11    32'h0000023b
`define DDRMC__SEQ_INIT_CNTRL11_SZ 10

`define DDRMC__SEQ_INIT_CNTRL12    32'h0000023c
`define DDRMC__SEQ_INIT_CNTRL12_SZ 10

`define DDRMC__SEQ_INIT_CNTRL13    32'h0000023d
`define DDRMC__SEQ_INIT_CNTRL13_SZ 10

`define DDRMC__SEQ_INIT_CNTRL14    32'h0000023e
`define DDRMC__SEQ_INIT_CNTRL14_SZ 10

`define DDRMC__SEQ_INIT_CNTRL15    32'h0000023f
`define DDRMC__SEQ_INIT_CNTRL15_SZ 10

`define DDRMC__SEQ_INIT_CNTRL16    32'h00000240
`define DDRMC__SEQ_INIT_CNTRL16_SZ 10

`define DDRMC__SEQ_INIT_CNTRL17    32'h00000241
`define DDRMC__SEQ_INIT_CNTRL17_SZ 10

`define DDRMC__SEQ_INIT_CNTRL18    32'h00000242
`define DDRMC__SEQ_INIT_CNTRL18_SZ 10

`define DDRMC__SEQ_INIT_CNTRL19    32'h00000243
`define DDRMC__SEQ_INIT_CNTRL19_SZ 10

`define DDRMC__SEQ_INIT_CNTRL2    32'h00000244
`define DDRMC__SEQ_INIT_CNTRL2_SZ 10

`define DDRMC__SEQ_INIT_CNTRL20    32'h00000245
`define DDRMC__SEQ_INIT_CNTRL20_SZ 10

`define DDRMC__SEQ_INIT_CNTRL21    32'h00000246
`define DDRMC__SEQ_INIT_CNTRL21_SZ 10

`define DDRMC__SEQ_INIT_CNTRL22    32'h00000247
`define DDRMC__SEQ_INIT_CNTRL22_SZ 10

`define DDRMC__SEQ_INIT_CNTRL23    32'h00000248
`define DDRMC__SEQ_INIT_CNTRL23_SZ 10

`define DDRMC__SEQ_INIT_CNTRL24    32'h00000249
`define DDRMC__SEQ_INIT_CNTRL24_SZ 10

`define DDRMC__SEQ_INIT_CNTRL25    32'h0000024a
`define DDRMC__SEQ_INIT_CNTRL25_SZ 10

`define DDRMC__SEQ_INIT_CNTRL26    32'h0000024b
`define DDRMC__SEQ_INIT_CNTRL26_SZ 10

`define DDRMC__SEQ_INIT_CNTRL27    32'h0000024c
`define DDRMC__SEQ_INIT_CNTRL27_SZ 10

`define DDRMC__SEQ_INIT_CNTRL28    32'h0000024d
`define DDRMC__SEQ_INIT_CNTRL28_SZ 10

`define DDRMC__SEQ_INIT_CNTRL29    32'h0000024e
`define DDRMC__SEQ_INIT_CNTRL29_SZ 10

`define DDRMC__SEQ_INIT_CNTRL3    32'h0000024f
`define DDRMC__SEQ_INIT_CNTRL3_SZ 10

`define DDRMC__SEQ_INIT_CNTRL30    32'h00000250
`define DDRMC__SEQ_INIT_CNTRL30_SZ 10

`define DDRMC__SEQ_INIT_CNTRL31    32'h00000251
`define DDRMC__SEQ_INIT_CNTRL31_SZ 10

`define DDRMC__SEQ_INIT_CNTRL32    32'h00000252
`define DDRMC__SEQ_INIT_CNTRL32_SZ 10

`define DDRMC__SEQ_INIT_CNTRL33    32'h00000253
`define DDRMC__SEQ_INIT_CNTRL33_SZ 10

`define DDRMC__SEQ_INIT_CNTRL34    32'h00000254
`define DDRMC__SEQ_INIT_CNTRL34_SZ 10

`define DDRMC__SEQ_INIT_CNTRL35    32'h00000255
`define DDRMC__SEQ_INIT_CNTRL35_SZ 10

`define DDRMC__SEQ_INIT_CNTRL36    32'h00000256
`define DDRMC__SEQ_INIT_CNTRL36_SZ 10

`define DDRMC__SEQ_INIT_CNTRL37    32'h00000257
`define DDRMC__SEQ_INIT_CNTRL37_SZ 10

`define DDRMC__SEQ_INIT_CNTRL38    32'h00000258
`define DDRMC__SEQ_INIT_CNTRL38_SZ 10

`define DDRMC__SEQ_INIT_CNTRL39    32'h00000259
`define DDRMC__SEQ_INIT_CNTRL39_SZ 10

`define DDRMC__SEQ_INIT_CNTRL4    32'h0000025a
`define DDRMC__SEQ_INIT_CNTRL4_SZ 10

`define DDRMC__SEQ_INIT_CNTRL40    32'h0000025b
`define DDRMC__SEQ_INIT_CNTRL40_SZ 10

`define DDRMC__SEQ_INIT_CNTRL41    32'h0000025c
`define DDRMC__SEQ_INIT_CNTRL41_SZ 10

`define DDRMC__SEQ_INIT_CNTRL42    32'h0000025d
`define DDRMC__SEQ_INIT_CNTRL42_SZ 10

`define DDRMC__SEQ_INIT_CNTRL43    32'h0000025e
`define DDRMC__SEQ_INIT_CNTRL43_SZ 10

`define DDRMC__SEQ_INIT_CNTRL44    32'h0000025f
`define DDRMC__SEQ_INIT_CNTRL44_SZ 10

`define DDRMC__SEQ_INIT_CNTRL45    32'h00000260
`define DDRMC__SEQ_INIT_CNTRL45_SZ 10

`define DDRMC__SEQ_INIT_CNTRL46    32'h00000261
`define DDRMC__SEQ_INIT_CNTRL46_SZ 10

`define DDRMC__SEQ_INIT_CNTRL47    32'h00000262
`define DDRMC__SEQ_INIT_CNTRL47_SZ 10

`define DDRMC__SEQ_INIT_CNTRL48    32'h00000263
`define DDRMC__SEQ_INIT_CNTRL48_SZ 10

`define DDRMC__SEQ_INIT_CNTRL49    32'h00000264
`define DDRMC__SEQ_INIT_CNTRL49_SZ 10

`define DDRMC__SEQ_INIT_CNTRL5    32'h00000265
`define DDRMC__SEQ_INIT_CNTRL5_SZ 10

`define DDRMC__SEQ_INIT_CNTRL50    32'h00000266
`define DDRMC__SEQ_INIT_CNTRL50_SZ 10

`define DDRMC__SEQ_INIT_CNTRL51    32'h00000267
`define DDRMC__SEQ_INIT_CNTRL51_SZ 10

`define DDRMC__SEQ_INIT_CNTRL52    32'h00000268
`define DDRMC__SEQ_INIT_CNTRL52_SZ 10

`define DDRMC__SEQ_INIT_CNTRL53    32'h00000269
`define DDRMC__SEQ_INIT_CNTRL53_SZ 10

`define DDRMC__SEQ_INIT_CNTRL54    32'h0000026a
`define DDRMC__SEQ_INIT_CNTRL54_SZ 10

`define DDRMC__SEQ_INIT_CNTRL55    32'h0000026b
`define DDRMC__SEQ_INIT_CNTRL55_SZ 10

`define DDRMC__SEQ_INIT_CNTRL56    32'h0000026c
`define DDRMC__SEQ_INIT_CNTRL56_SZ 10

`define DDRMC__SEQ_INIT_CNTRL57    32'h0000026d
`define DDRMC__SEQ_INIT_CNTRL57_SZ 10

`define DDRMC__SEQ_INIT_CNTRL58    32'h0000026e
`define DDRMC__SEQ_INIT_CNTRL58_SZ 10

`define DDRMC__SEQ_INIT_CNTRL59    32'h0000026f
`define DDRMC__SEQ_INIT_CNTRL59_SZ 10

`define DDRMC__SEQ_INIT_CNTRL6    32'h00000270
`define DDRMC__SEQ_INIT_CNTRL6_SZ 10

`define DDRMC__SEQ_INIT_CNTRL60    32'h00000271
`define DDRMC__SEQ_INIT_CNTRL60_SZ 10

`define DDRMC__SEQ_INIT_CNTRL61    32'h00000272
`define DDRMC__SEQ_INIT_CNTRL61_SZ 10

`define DDRMC__SEQ_INIT_CNTRL62    32'h00000273
`define DDRMC__SEQ_INIT_CNTRL62_SZ 10

`define DDRMC__SEQ_INIT_CNTRL63    32'h00000274
`define DDRMC__SEQ_INIT_CNTRL63_SZ 10

`define DDRMC__SEQ_INIT_CNTRL64    32'h00000275
`define DDRMC__SEQ_INIT_CNTRL64_SZ 10

`define DDRMC__SEQ_INIT_CNTRL65    32'h00000276
`define DDRMC__SEQ_INIT_CNTRL65_SZ 10

`define DDRMC__SEQ_INIT_CNTRL66    32'h00000277
`define DDRMC__SEQ_INIT_CNTRL66_SZ 10

`define DDRMC__SEQ_INIT_CNTRL67    32'h00000278
`define DDRMC__SEQ_INIT_CNTRL67_SZ 10

`define DDRMC__SEQ_INIT_CNTRL68    32'h00000279
`define DDRMC__SEQ_INIT_CNTRL68_SZ 10

`define DDRMC__SEQ_INIT_CNTRL69    32'h0000027a
`define DDRMC__SEQ_INIT_CNTRL69_SZ 10

`define DDRMC__SEQ_INIT_CNTRL7    32'h0000027b
`define DDRMC__SEQ_INIT_CNTRL7_SZ 10

`define DDRMC__SEQ_INIT_CNTRL70    32'h0000027c
`define DDRMC__SEQ_INIT_CNTRL70_SZ 10

`define DDRMC__SEQ_INIT_CNTRL71    32'h0000027d
`define DDRMC__SEQ_INIT_CNTRL71_SZ 10

`define DDRMC__SEQ_INIT_CNTRL72    32'h0000027e
`define DDRMC__SEQ_INIT_CNTRL72_SZ 10

`define DDRMC__SEQ_INIT_CNTRL73    32'h0000027f
`define DDRMC__SEQ_INIT_CNTRL73_SZ 10

`define DDRMC__SEQ_INIT_CNTRL74    32'h00000280
`define DDRMC__SEQ_INIT_CNTRL74_SZ 10

`define DDRMC__SEQ_INIT_CNTRL75    32'h00000281
`define DDRMC__SEQ_INIT_CNTRL75_SZ 10

`define DDRMC__SEQ_INIT_CNTRL76    32'h00000282
`define DDRMC__SEQ_INIT_CNTRL76_SZ 10

`define DDRMC__SEQ_INIT_CNTRL77    32'h00000283
`define DDRMC__SEQ_INIT_CNTRL77_SZ 10

`define DDRMC__SEQ_INIT_CNTRL78    32'h00000284
`define DDRMC__SEQ_INIT_CNTRL78_SZ 10

`define DDRMC__SEQ_INIT_CNTRL79    32'h00000285
`define DDRMC__SEQ_INIT_CNTRL79_SZ 10

`define DDRMC__SEQ_INIT_CNTRL8    32'h00000286
`define DDRMC__SEQ_INIT_CNTRL8_SZ 10

`define DDRMC__SEQ_INIT_CNTRL80    32'h00000287
`define DDRMC__SEQ_INIT_CNTRL80_SZ 10

`define DDRMC__SEQ_INIT_CNTRL81    32'h00000288
`define DDRMC__SEQ_INIT_CNTRL81_SZ 10

`define DDRMC__SEQ_INIT_CNTRL82    32'h00000289
`define DDRMC__SEQ_INIT_CNTRL82_SZ 10

`define DDRMC__SEQ_INIT_CNTRL83    32'h0000028a
`define DDRMC__SEQ_INIT_CNTRL83_SZ 10

`define DDRMC__SEQ_INIT_CNTRL84    32'h0000028b
`define DDRMC__SEQ_INIT_CNTRL84_SZ 10

`define DDRMC__SEQ_INIT_CNTRL85    32'h0000028c
`define DDRMC__SEQ_INIT_CNTRL85_SZ 10

`define DDRMC__SEQ_INIT_CNTRL86    32'h0000028d
`define DDRMC__SEQ_INIT_CNTRL86_SZ 10

`define DDRMC__SEQ_INIT_CNTRL87    32'h0000028e
`define DDRMC__SEQ_INIT_CNTRL87_SZ 10

`define DDRMC__SEQ_INIT_CNTRL88    32'h0000028f
`define DDRMC__SEQ_INIT_CNTRL88_SZ 10

`define DDRMC__SEQ_INIT_CNTRL89    32'h00000290
`define DDRMC__SEQ_INIT_CNTRL89_SZ 10

`define DDRMC__SEQ_INIT_CNTRL9    32'h00000291
`define DDRMC__SEQ_INIT_CNTRL9_SZ 10

`define DDRMC__SEQ_INIT_CNTRL90    32'h00000292
`define DDRMC__SEQ_INIT_CNTRL90_SZ 10

`define DDRMC__SEQ_INIT_CNTRL91    32'h00000293
`define DDRMC__SEQ_INIT_CNTRL91_SZ 10

`define DDRMC__SEQ_INIT_CNTRL92    32'h00000294
`define DDRMC__SEQ_INIT_CNTRL92_SZ 10

`define DDRMC__SEQ_INIT_CNTRL93    32'h00000295
`define DDRMC__SEQ_INIT_CNTRL93_SZ 10

`define DDRMC__SEQ_INIT_CNTRL94    32'h00000296
`define DDRMC__SEQ_INIT_CNTRL94_SZ 10

`define DDRMC__SEQ_INIT_CNTRL95    32'h00000297
`define DDRMC__SEQ_INIT_CNTRL95_SZ 10

`define DDRMC__SEQ_INIT_CNTRL96    32'h00000298
`define DDRMC__SEQ_INIT_CNTRL96_SZ 10

`define DDRMC__SEQ_INIT_CNTRL97    32'h00000299
`define DDRMC__SEQ_INIT_CNTRL97_SZ 10

`define DDRMC__SEQ_INIT_CNTRL98    32'h0000029a
`define DDRMC__SEQ_INIT_CNTRL98_SZ 10

`define DDRMC__SEQ_INIT_CNTRL99    32'h0000029b
`define DDRMC__SEQ_INIT_CNTRL99_SZ 10

`define DDRMC__SEQ_INIT_CONFIG    32'h0000029c
`define DDRMC__SEQ_INIT_CONFIG_SZ 17

`define DDRMC__SEQ_MODE    32'h0000029d
`define DDRMC__SEQ_MODE_SZ 3

`define DDRMC__TXNQ_RD_PRIORITY    32'h0000029e
`define DDRMC__TXNQ_RD_PRIORITY_SZ 26

`define DDRMC__TXNQ_WR_PRIORITY    32'h0000029f
`define DDRMC__TXNQ_WR_PRIORITY_SZ 25

`define DDRMC__T_TXBIT    32'h000002a0
`define DDRMC__T_TXBIT_SZ 1

`define DDRMC__UB_CLK_MUX    32'h000002a1
`define DDRMC__UB_CLK_MUX_SZ 2

`define DDRMC__WRITE_BANDWIDTH    32'h000002a2
`define DDRMC__WRITE_BANDWIDTH_SZ 64

`define DDRMC__XMPU_CONFIG0    32'h000002a3
`define DDRMC__XMPU_CONFIG0_SZ 5

`define DDRMC__XMPU_CONFIG1    32'h000002a4
`define DDRMC__XMPU_CONFIG1_SZ 5

`define DDRMC__XMPU_CONFIG10    32'h000002a5
`define DDRMC__XMPU_CONFIG10_SZ 5

`define DDRMC__XMPU_CONFIG11    32'h000002a6
`define DDRMC__XMPU_CONFIG11_SZ 5

`define DDRMC__XMPU_CONFIG12    32'h000002a7
`define DDRMC__XMPU_CONFIG12_SZ 5

`define DDRMC__XMPU_CONFIG13    32'h000002a8
`define DDRMC__XMPU_CONFIG13_SZ 5

`define DDRMC__XMPU_CONFIG14    32'h000002a9
`define DDRMC__XMPU_CONFIG14_SZ 5

`define DDRMC__XMPU_CONFIG15    32'h000002aa
`define DDRMC__XMPU_CONFIG15_SZ 5

`define DDRMC__XMPU_CONFIG2    32'h000002ab
`define DDRMC__XMPU_CONFIG2_SZ 5

`define DDRMC__XMPU_CONFIG3    32'h000002ac
`define DDRMC__XMPU_CONFIG3_SZ 5

`define DDRMC__XMPU_CONFIG4    32'h000002ad
`define DDRMC__XMPU_CONFIG4_SZ 5

`define DDRMC__XMPU_CONFIG5    32'h000002ae
`define DDRMC__XMPU_CONFIG5_SZ 5

`define DDRMC__XMPU_CONFIG6    32'h000002af
`define DDRMC__XMPU_CONFIG6_SZ 5

`define DDRMC__XMPU_CONFIG7    32'h000002b0
`define DDRMC__XMPU_CONFIG7_SZ 5

`define DDRMC__XMPU_CONFIG8    32'h000002b1
`define DDRMC__XMPU_CONFIG8_SZ 5

`define DDRMC__XMPU_CONFIG9    32'h000002b2
`define DDRMC__XMPU_CONFIG9_SZ 5

`define DDRMC__XMPU_CTRL    32'h000002b3
`define DDRMC__XMPU_CTRL_SZ 4

`define DDRMC__XMPU_END_HI0    32'h000002b4
`define DDRMC__XMPU_END_HI0_SZ 16

`define DDRMC__XMPU_END_HI1    32'h000002b5
`define DDRMC__XMPU_END_HI1_SZ 16

`define DDRMC__XMPU_END_HI10    32'h000002b6
`define DDRMC__XMPU_END_HI10_SZ 16

`define DDRMC__XMPU_END_HI11    32'h000002b7
`define DDRMC__XMPU_END_HI11_SZ 16

`define DDRMC__XMPU_END_HI12    32'h000002b8
`define DDRMC__XMPU_END_HI12_SZ 16

`define DDRMC__XMPU_END_HI13    32'h000002b9
`define DDRMC__XMPU_END_HI13_SZ 16

`define DDRMC__XMPU_END_HI14    32'h000002ba
`define DDRMC__XMPU_END_HI14_SZ 16

`define DDRMC__XMPU_END_HI15    32'h000002bb
`define DDRMC__XMPU_END_HI15_SZ 16

`define DDRMC__XMPU_END_HI2    32'h000002bc
`define DDRMC__XMPU_END_HI2_SZ 16

`define DDRMC__XMPU_END_HI3    32'h000002bd
`define DDRMC__XMPU_END_HI3_SZ 16

`define DDRMC__XMPU_END_HI4    32'h000002be
`define DDRMC__XMPU_END_HI4_SZ 16

`define DDRMC__XMPU_END_HI5    32'h000002bf
`define DDRMC__XMPU_END_HI5_SZ 16

`define DDRMC__XMPU_END_HI6    32'h000002c0
`define DDRMC__XMPU_END_HI6_SZ 16

`define DDRMC__XMPU_END_HI7    32'h000002c1
`define DDRMC__XMPU_END_HI7_SZ 16

`define DDRMC__XMPU_END_HI8    32'h000002c2
`define DDRMC__XMPU_END_HI8_SZ 16

`define DDRMC__XMPU_END_HI9    32'h000002c3
`define DDRMC__XMPU_END_HI9_SZ 16

`define DDRMC__XMPU_END_LO0    32'h000002c4
`define DDRMC__XMPU_END_LO0_SZ 32

`define DDRMC__XMPU_END_LO1    32'h000002c5
`define DDRMC__XMPU_END_LO1_SZ 32

`define DDRMC__XMPU_END_LO10    32'h000002c6
`define DDRMC__XMPU_END_LO10_SZ 32

`define DDRMC__XMPU_END_LO11    32'h000002c7
`define DDRMC__XMPU_END_LO11_SZ 32

`define DDRMC__XMPU_END_LO12    32'h000002c8
`define DDRMC__XMPU_END_LO12_SZ 32

`define DDRMC__XMPU_END_LO13    32'h000002c9
`define DDRMC__XMPU_END_LO13_SZ 32

`define DDRMC__XMPU_END_LO14    32'h000002ca
`define DDRMC__XMPU_END_LO14_SZ 32

`define DDRMC__XMPU_END_LO15    32'h000002cb
`define DDRMC__XMPU_END_LO15_SZ 32

`define DDRMC__XMPU_END_LO2    32'h000002cc
`define DDRMC__XMPU_END_LO2_SZ 32

`define DDRMC__XMPU_END_LO3    32'h000002cd
`define DDRMC__XMPU_END_LO3_SZ 32

`define DDRMC__XMPU_END_LO4    32'h000002ce
`define DDRMC__XMPU_END_LO4_SZ 32

`define DDRMC__XMPU_END_LO5    32'h000002cf
`define DDRMC__XMPU_END_LO5_SZ 32

`define DDRMC__XMPU_END_LO6    32'h000002d0
`define DDRMC__XMPU_END_LO6_SZ 32

`define DDRMC__XMPU_END_LO7    32'h000002d1
`define DDRMC__XMPU_END_LO7_SZ 32

`define DDRMC__XMPU_END_LO8    32'h000002d2
`define DDRMC__XMPU_END_LO8_SZ 32

`define DDRMC__XMPU_END_LO9    32'h000002d3
`define DDRMC__XMPU_END_LO9_SZ 32

`define DDRMC__XMPU_MASTER0    32'h000002d4
`define DDRMC__XMPU_MASTER0_SZ 26

`define DDRMC__XMPU_MASTER1    32'h000002d5
`define DDRMC__XMPU_MASTER1_SZ 26

`define DDRMC__XMPU_MASTER10    32'h000002d6
`define DDRMC__XMPU_MASTER10_SZ 26

`define DDRMC__XMPU_MASTER11    32'h000002d7
`define DDRMC__XMPU_MASTER11_SZ 26

`define DDRMC__XMPU_MASTER12    32'h000002d8
`define DDRMC__XMPU_MASTER12_SZ 26

`define DDRMC__XMPU_MASTER13    32'h000002d9
`define DDRMC__XMPU_MASTER13_SZ 26

`define DDRMC__XMPU_MASTER14    32'h000002da
`define DDRMC__XMPU_MASTER14_SZ 26

`define DDRMC__XMPU_MASTER15    32'h000002db
`define DDRMC__XMPU_MASTER15_SZ 26

`define DDRMC__XMPU_MASTER2    32'h000002dc
`define DDRMC__XMPU_MASTER2_SZ 26

`define DDRMC__XMPU_MASTER3    32'h000002dd
`define DDRMC__XMPU_MASTER3_SZ 26

`define DDRMC__XMPU_MASTER4    32'h000002de
`define DDRMC__XMPU_MASTER4_SZ 26

`define DDRMC__XMPU_MASTER5    32'h000002df
`define DDRMC__XMPU_MASTER5_SZ 26

`define DDRMC__XMPU_MASTER6    32'h000002e0
`define DDRMC__XMPU_MASTER6_SZ 26

`define DDRMC__XMPU_MASTER7    32'h000002e1
`define DDRMC__XMPU_MASTER7_SZ 26

`define DDRMC__XMPU_MASTER8    32'h000002e2
`define DDRMC__XMPU_MASTER8_SZ 26

`define DDRMC__XMPU_MASTER9    32'h000002e3
`define DDRMC__XMPU_MASTER9_SZ 26

`define DDRMC__XMPU_START_HI0    32'h000002e4
`define DDRMC__XMPU_START_HI0_SZ 16

`define DDRMC__XMPU_START_HI1    32'h000002e5
`define DDRMC__XMPU_START_HI1_SZ 16

`define DDRMC__XMPU_START_HI10    32'h000002e6
`define DDRMC__XMPU_START_HI10_SZ 16

`define DDRMC__XMPU_START_HI11    32'h000002e7
`define DDRMC__XMPU_START_HI11_SZ 16

`define DDRMC__XMPU_START_HI12    32'h000002e8
`define DDRMC__XMPU_START_HI12_SZ 16

`define DDRMC__XMPU_START_HI13    32'h000002e9
`define DDRMC__XMPU_START_HI13_SZ 16

`define DDRMC__XMPU_START_HI14    32'h000002ea
`define DDRMC__XMPU_START_HI14_SZ 16

`define DDRMC__XMPU_START_HI15    32'h000002eb
`define DDRMC__XMPU_START_HI15_SZ 16

`define DDRMC__XMPU_START_HI2    32'h000002ec
`define DDRMC__XMPU_START_HI2_SZ 16

`define DDRMC__XMPU_START_HI3    32'h000002ed
`define DDRMC__XMPU_START_HI3_SZ 16

`define DDRMC__XMPU_START_HI4    32'h000002ee
`define DDRMC__XMPU_START_HI4_SZ 16

`define DDRMC__XMPU_START_HI5    32'h000002ef
`define DDRMC__XMPU_START_HI5_SZ 16

`define DDRMC__XMPU_START_HI6    32'h000002f0
`define DDRMC__XMPU_START_HI6_SZ 16

`define DDRMC__XMPU_START_HI7    32'h000002f1
`define DDRMC__XMPU_START_HI7_SZ 16

`define DDRMC__XMPU_START_HI8    32'h000002f2
`define DDRMC__XMPU_START_HI8_SZ 16

`define DDRMC__XMPU_START_HI9    32'h000002f3
`define DDRMC__XMPU_START_HI9_SZ 16

`define DDRMC__XMPU_START_LO0    32'h000002f4
`define DDRMC__XMPU_START_LO0_SZ 32

`define DDRMC__XMPU_START_LO1    32'h000002f5
`define DDRMC__XMPU_START_LO1_SZ 32

`define DDRMC__XMPU_START_LO10    32'h000002f6
`define DDRMC__XMPU_START_LO10_SZ 32

`define DDRMC__XMPU_START_LO11    32'h000002f7
`define DDRMC__XMPU_START_LO11_SZ 32

`define DDRMC__XMPU_START_LO12    32'h000002f8
`define DDRMC__XMPU_START_LO12_SZ 32

`define DDRMC__XMPU_START_LO13    32'h000002f9
`define DDRMC__XMPU_START_LO13_SZ 32

`define DDRMC__XMPU_START_LO14    32'h000002fa
`define DDRMC__XMPU_START_LO14_SZ 32

`define DDRMC__XMPU_START_LO15    32'h000002fb
`define DDRMC__XMPU_START_LO15_SZ 32

`define DDRMC__XMPU_START_LO2    32'h000002fc
`define DDRMC__XMPU_START_LO2_SZ 32

`define DDRMC__XMPU_START_LO3    32'h000002fd
`define DDRMC__XMPU_START_LO3_SZ 32

`define DDRMC__XMPU_START_LO4    32'h000002fe
`define DDRMC__XMPU_START_LO4_SZ 32

`define DDRMC__XMPU_START_LO5    32'h000002ff
`define DDRMC__XMPU_START_LO5_SZ 32

`define DDRMC__XMPU_START_LO6    32'h00000300
`define DDRMC__XMPU_START_LO6_SZ 32

`define DDRMC__XMPU_START_LO7    32'h00000301
`define DDRMC__XMPU_START_LO7_SZ 32

`define DDRMC__XMPU_START_LO8    32'h00000302
`define DDRMC__XMPU_START_LO8_SZ 32

`define DDRMC__XMPU_START_LO9    32'h00000303
`define DDRMC__XMPU_START_LO9_SZ 32

`define DDRMC__XPI_DATA_NIB_CHAN    32'h00000304
`define DDRMC__XPI_DATA_NIB_CHAN_SZ 18

`define DDRMC__XPI_DQS    32'h00000305
`define DDRMC__XPI_DQS_SZ 8

`define DDRMC__XPI_NIB_CHAN    32'h00000306
`define DDRMC__XPI_NIB_CHAN_SZ 27

`define DDRMC__XPI_OE    32'h00000307
`define DDRMC__XPI_OE_SZ 16

`define DDRMC__XPI_OE_ALL_NIB    32'h00000308
`define DDRMC__XPI_OE_ALL_NIB_SZ 11

`define DDRMC__XPI_PMI_CONFIG    32'h00000309
`define DDRMC__XPI_PMI_CONFIG_SZ 9

`define DDRMC__XPI_READ_DBI    32'h0000030a
`define DDRMC__XPI_READ_DBI_SZ 2

`define DDRMC__XPI_READ_OFFSET    32'h0000030b
`define DDRMC__XPI_READ_OFFSET_SZ 14

`define DDRMC__XPI_WRDATA_ALL_NIB    32'h0000030c
`define DDRMC__XPI_WRDATA_ALL_NIB_SZ 11

`define DDRMC__XPI_WRITE_DM_DBI    32'h0000030d
`define DDRMC__XPI_WRITE_DM_DBI_SZ 4

`endif  // B_DDRMC_DEFINES_VH