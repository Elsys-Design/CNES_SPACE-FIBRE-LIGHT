localparam A_CFG0 = 'd1856;
localparam A_CFG1 = 'd1316376142;
localparam A_CFG2 = 'd3758096384;
localparam A_CFG3 = 'd3758096384;
localparam A_CFG4 = 'd1610612736;
localparam A_CFG5 = 'd3758096384;
localparam CH0_ADAPT_APT_CFG = 'd0;
localparam CH0_ADAPT_CAL_CFG = 'd2179884032;
localparam CH0_ADAPT_DFE_CFG = 'd64;
localparam CH0_ADAPT_GC_CFG0 = 'd9441392;
localparam CH0_ADAPT_GC_CFG1 = 'd178259936;
localparam CH0_ADAPT_GC_CFG2 = 'd2097384;
localparam CH0_ADAPT_GC_CFG3 = 'd178258912;
localparam CH0_ADAPT_GEN_CFG0 = 'd1179648;
localparam CH0_ADAPT_GEN_CFG1 = 'd0;
localparam CH0_ADAPT_GEN_CFG2 = 'd2281701375;
localparam CH0_ADAPT_GEN_CFG3 = 'd268435456;
localparam CH0_ADAPT_H01_CFG = 'd18875040;
localparam CH0_ADAPT_H23_CFG = 'd27263392;
localparam CH0_ADAPT_H45_CFG = 'd27263392;
localparam CH0_ADAPT_H67_CFG = 'd27263392;
localparam CH0_ADAPT_H89_CFG = 'd27263392;
localparam CH0_ADAPT_HAB_CFG = 'd27263392;
localparam CH0_ADAPT_HCD_CFG = 'd27263392;
localparam CH0_ADAPT_HEF_CFG = 'd27263904;
localparam CH0_ADAPT_KH_CFG0 = 'd537426239;
localparam CH0_ADAPT_KH_CFG1 = 'd0;
localparam CH0_ADAPT_KH_CFG2 = 'd17312;
localparam CH0_ADAPT_KH_CFG3 = 'd0;
localparam CH0_ADAPT_KH_CFG4 = 'd31648;
localparam CH0_ADAPT_KH_CFG5 = 'd0;
localparam CH0_ADAPT_KL_CFG0 = 'd32928;
localparam CH0_ADAPT_KL_CFG1 = 'd17312;
localparam CH0_ADAPT_LCK_CFG0 = 'd16384;
localparam CH0_ADAPT_LCK_CFG1 = 'd16384;
localparam CH0_ADAPT_LCK_CFG2 = 'd0;
localparam CH0_ADAPT_LCK_CFG3 = 'd0;
localparam CH0_ADAPT_LOP_CFG = 'd3992979040;
localparam CH0_ADAPT_OS_CFG = 'd2147483936;
localparam CH0_CHCLK_ILO_CFG = 'd6553651;
localparam CH0_CHCLK_MISC_CFG = 'd4169260831;
localparam CH0_CHCLK_RSV_CFG = 'd0;
localparam CH0_CHCLK_RXCAL_CFG = 'd138166272;
localparam CH0_CHCLK_RXCAL_CFG1 = 'd0;
localparam CH0_CHCLK_RXCAL_CFG2 = 'd0;
localparam CH0_CHCLK_RXPI_CFG = 'd5244972;
localparam CH0_CHCLK_TXCAL_CFG = 'd4194336;
localparam CH0_CHCLK_TXPI_CFG0 = 'd4655151;
localparam CH0_CHL_RSV_CFG0 = 'd3330277385;
localparam CH0_CHL_RSV_CFG1 = 'd1560;
localparam CH0_CHL_RSV_CFG2 = 'd6227344;
localparam CH0_CHL_RSV_CFG3 = 'd0;
localparam CH0_CHL_RSV_CFG4 = 'd0;
localparam CH0_DA_CFG = 'd655370;
localparam CH0_EYESCAN_CFG0 = 'd2048;
localparam CH0_EYESCAN_CFG1 = 'd0;
localparam CH0_EYESCAN_CFG10 = 'd0;
localparam CH0_EYESCAN_CFG11 = 'd0;
localparam CH0_EYESCAN_CFG12 = 'd0;
localparam CH0_EYESCAN_CFG13 = 'd0;
localparam CH0_EYESCAN_CFG14 = 'd0;
localparam CH0_EYESCAN_CFG15 = 'd0;
localparam CH0_EYESCAN_CFG16 = 'd0;
localparam CH0_EYESCAN_CFG2 = 'd0;
localparam CH0_EYESCAN_CFG3 = 'd0;
localparam CH0_EYESCAN_CFG4 = 'd0;
localparam CH0_EYESCAN_CFG5 = 'd0;
localparam CH0_EYESCAN_CFG6 = 'd0;
localparam CH0_EYESCAN_CFG7 = 'd0;
localparam CH0_EYESCAN_CFG8 = 'd0;
localparam CH0_EYESCAN_CFG9 = 'd0;
localparam CH0_FABRIC_INTF_CFG0 = 'd4273993723;
localparam CH0_FABRIC_INTF_CFG1 = 'd197632;
localparam CH0_FABRIC_INTF_CFG2 = 'd537919472;
localparam CH0_FABRIC_INTF_CFG3 = 'd786432;
localparam CH0_FABRIC_INTF_CFG4 = 'd20480;
localparam CH0_FABRIC_INTF_CFG5 = 'd25602;
localparam CH0_INSTANTIATED = 'd0;
localparam CH0_MONITOR_CFG = 'd0;
localparam CH0_PIPE_CTRL_CFG0 = 'd262240;
localparam CH0_PIPE_CTRL_CFG1 = 'd2097811;
localparam CH0_PIPE_CTRL_CFG10 = 'd85983215;
localparam CH0_PIPE_CTRL_CFG2 = 'd9950092;
localparam CH0_PIPE_CTRL_CFG3 = 'd1573167;
localparam CH0_PIPE_CTRL_CFG4 = 'd1078198272;
localparam CH0_PIPE_CTRL_CFG5 = 'd2684354560;
localparam CH0_PIPE_CTRL_CFG6 = 'd1007681636;
localparam CH0_PIPE_CTRL_CFG7 = 'd67149834;
localparam CH0_PIPE_CTRL_CFG8 = 'd33554432;
localparam CH0_PIPE_CTRL_CFG9 = 'd0;
localparam CH0_PIPE_TX_EQ_CFG0 = 'd175467487;
localparam CH0_PIPE_TX_EQ_CFG1 = 'd152233553;
localparam CH0_PIPE_TX_EQ_CFG2 = 'd8258;
localparam CH0_PIPE_TX_EQ_CFG3 = 'd393618;
localparam CH0_RESET_BYP_HDSHK_CFG = 'd0;
localparam CH0_RESET_CFG = 'd135266341;
localparam CH0_RESET_LOOPER_ID_CFG = 'd2113632;
localparam CH0_RESET_LOOP_ID_CFG0 = 'd528;
localparam CH0_RESET_LOOP_ID_CFG1 = 'd106181136;
localparam CH0_RESET_LOOP_ID_CFG2 = 'd17185;
localparam CH0_RESET_TIME_CFG0 = 'd34636801;
localparam CH0_RESET_TIME_CFG1 = 'd34636833;
localparam CH0_RESET_TIME_CFG2 = 'd34636833;
localparam CH0_RESET_TIME_CFG3 = 'd2231903265;
localparam CH0_RXOUTCLK_FREQ = 390.625;
localparam CH0_RXOUTCLK_REF_FREQ = 125;
localparam CH0_RXOUTCLK_REF_SOURCE = "HSCLK0_LCPLLGTREFCLK0";
localparam CH0_RX_CDR_CFG0 = 'd3019898946;
localparam CH0_RX_CDR_CFG1 = 'd1610612992;
localparam CH0_RX_CDR_CFG2 = 'd134236777;
localparam CH0_RX_CDR_CFG3 = 'd744694;
localparam CH0_RX_CDR_CFG4 = 'd607924224;
localparam CH0_RX_CRC_CFG0 = 'd30848;
localparam CH0_RX_CRC_CFG1 = 'd505290270;
localparam CH0_RX_CRC_CFG2 = 'd505290270;
localparam CH0_RX_CRC_CFG3 = 'd4294967295;
localparam CH0_RX_CTLE_CFG0 = 'd31195392;
localparam CH0_RX_CTLE_CFG1 = 'd1073741824;
localparam CH0_RX_DACI2V_CFG0 = 'd67145418;
localparam CH0_RX_DFE_CFG0 = 'd3489813512;
localparam CH0_RX_ELASTIC_BUF_CFG0 = 'd2155632704;
localparam CH0_RX_ELASTIC_BUF_CFG1 = 'd2;
localparam CH0_RX_ELASTIC_BUF_CFG2 = 'd0;
localparam CH0_RX_ELASTIC_BUF_CFG3 = 'd2682257408;
localparam CH0_RX_ELASTIC_BUF_CFG4 = 'd0;
localparam CH0_RX_ELASTIC_BUF_CFG5 = 'd0;
localparam CH0_RX_ELASTIC_BUF_CFG6 = 'd4293918720;
localparam CH0_RX_ELASTIC_BUF_CFG7 = 'd67108869;
localparam CH0_RX_ELASTIC_BUF_CFG8 = 'd2033040;
localparam CH0_RX_ELASTIC_BUF_CFG9 = 'd2033040;
localparam CH0_RX_MISC_CFG0 = 'd1342177280;
localparam CH0_RX_OOB_CFG0 = 'd609534468;
localparam CH0_RX_OOB_CFG1 = 'd16925124;
localparam CH0_RX_PAD_CFG0 = 'd0;
localparam CH0_RX_PAD_CFG1 = 'd272910714;
localparam CH0_RX_PCS_CFG0 = 'd674623792;
localparam CH0_RX_PCS_CFG1 = 'd1812204543;
localparam CH0_RX_PCS_CFG2 = 'd1073742049;
localparam CH0_RX_PCS_CFG3 = 'd471666447;
localparam CH0_RX_PCS_CFG4 = 'd1115725826;
localparam CH0_RX_PHALIGN_CFG0 = 'd3;
localparam CH0_RX_PHALIGN_CFG1 = 'd8617984;
localparam CH0_RX_PHALIGN_CFG2 = 'd117248;
localparam CH0_RX_PHALIGN_CFG3 = 'd229376;
localparam CH0_RX_PHALIGN_CFG4 = 'd522;
localparam CH0_RX_PHALIGN_CFG5 = 'd50462720;
localparam CH0_TXOUTCLK_FREQ = 390.625;
localparam CH0_TXOUTCLK_REF_FREQ = 125;
localparam CH0_TXOUTCLK_REF_SOURCE = "HSCLK0_LCPLLGTREFCLK0";
localparam CH0_TX_10G_CFG0 = 'd0;
localparam CH0_TX_10G_CFG1 = 'd1073741824;
localparam CH0_TX_10G_CFG2 = 'd0;
localparam CH0_TX_10G_CFG3 = 'd0;
localparam CH0_TX_ANA_CFG0 = 'd208;
localparam CH0_TX_CRC_CFG0 = 'd30720;
localparam CH0_TX_CRC_CFG1 = 'd505290270;
localparam CH0_TX_CRC_CFG2 = 'd505290270;
localparam CH0_TX_CRC_CFG3 = 'd4294967295;
localparam CH0_TX_DRV_CFG0 = 'd4194304;
localparam CH0_TX_DRV_CFG1 = 'd6144;
localparam CH0_TX_PCS_CFG0 = 'd2187329825;
localparam CH0_TX_PCS_CFG1 = 'd674583932;
localparam CH0_TX_PCS_CFG2 = 'd357954218;
localparam CH0_TX_PCS_CFG3 = 'd1747587;
localparam CH0_TX_PHALIGN_CFG0 = 'd0;
localparam CH0_TX_PHALIGN_CFG1 = 'd290816;
localparam CH0_TX_PHALIGN_CFG2 = 'd229432;
localparam CH0_TX_PHALIGN_CFG3 = 'd0;
localparam CH0_TX_PHALIGN_CFG4 = 'd402653408;
localparam CH0_TX_PHALIGN_CFG5 = 'd128;
localparam CH0_TX_PIPPM_CFG = 'd33554432;
localparam CH0_TX_SER_CFG0 = 'd0;
localparam CH1_ADAPT_APT_CFG = 'd0;
localparam CH1_ADAPT_CAL_CFG = 'd2179884032;
localparam CH1_ADAPT_DFE_CFG = 'd64;
localparam CH1_ADAPT_GC_CFG0 = 'd9441392;
localparam CH1_ADAPT_GC_CFG1 = 'd178259936;
localparam CH1_ADAPT_GC_CFG2 = 'd2097384;
localparam CH1_ADAPT_GC_CFG3 = 'd178258912;
localparam CH1_ADAPT_GEN_CFG0 = 'd1179648;
localparam CH1_ADAPT_GEN_CFG1 = 'd0;
localparam CH1_ADAPT_GEN_CFG2 = 'd2281701375;
localparam CH1_ADAPT_GEN_CFG3 = 'd268435456;
localparam CH1_ADAPT_H01_CFG = 'd18875040;
localparam CH1_ADAPT_H23_CFG = 'd27263392;
localparam CH1_ADAPT_H45_CFG = 'd27263392;
localparam CH1_ADAPT_H67_CFG = 'd27263392;
localparam CH1_ADAPT_H89_CFG = 'd27263392;
localparam CH1_ADAPT_HAB_CFG = 'd27263392;
localparam CH1_ADAPT_HCD_CFG = 'd27263392;
localparam CH1_ADAPT_HEF_CFG = 'd27263904;
localparam CH1_ADAPT_KH_CFG0 = 'd537426239;
localparam CH1_ADAPT_KH_CFG1 = 'd0;
localparam CH1_ADAPT_KH_CFG2 = 'd17312;
localparam CH1_ADAPT_KH_CFG3 = 'd0;
localparam CH1_ADAPT_KH_CFG4 = 'd31648;
localparam CH1_ADAPT_KH_CFG5 = 'd0;
localparam CH1_ADAPT_KL_CFG0 = 'd32928;
localparam CH1_ADAPT_KL_CFG1 = 'd17312;
localparam CH1_ADAPT_LCK_CFG0 = 'd16384;
localparam CH1_ADAPT_LCK_CFG1 = 'd16384;
localparam CH1_ADAPT_LCK_CFG2 = 'd0;
localparam CH1_ADAPT_LCK_CFG3 = 'd0;
localparam CH1_ADAPT_LOP_CFG = 'd3992979040;
localparam CH1_ADAPT_OS_CFG = 'd2147483936;
localparam CH1_CHCLK_ILO_CFG = 'd6553651;
localparam CH1_CHCLK_MISC_CFG = 'd4169260831;
localparam CH1_CHCLK_RSV_CFG = 'd0;
localparam CH1_CHCLK_RXCAL_CFG = 'd138166272;
localparam CH1_CHCLK_RXCAL_CFG1 = 'd0;
localparam CH1_CHCLK_RXCAL_CFG2 = 'd0;
localparam CH1_CHCLK_RXPI_CFG = 'd5244972;
localparam CH1_CHCLK_TXCAL_CFG = 'd4194336;
localparam CH1_CHCLK_TXPI_CFG0 = 'd4655151;
localparam CH1_CHL_RSV_CFG0 = 'd3330277385;
localparam CH1_CHL_RSV_CFG1 = 'd1560;
localparam CH1_CHL_RSV_CFG2 = 'd6227344;
localparam CH1_CHL_RSV_CFG3 = 'd0;
localparam CH1_CHL_RSV_CFG4 = 'd0;
localparam CH1_DA_CFG = 'd655370;
localparam CH1_EYESCAN_CFG0 = 'd2048;
localparam CH1_EYESCAN_CFG1 = 'd0;
localparam CH1_EYESCAN_CFG10 = 'd0;
localparam CH1_EYESCAN_CFG11 = 'd0;
localparam CH1_EYESCAN_CFG12 = 'd0;
localparam CH1_EYESCAN_CFG13 = 'd0;
localparam CH1_EYESCAN_CFG14 = 'd0;
localparam CH1_EYESCAN_CFG15 = 'd0;
localparam CH1_EYESCAN_CFG16 = 'd0;
localparam CH1_EYESCAN_CFG2 = 'd0;
localparam CH1_EYESCAN_CFG3 = 'd0;
localparam CH1_EYESCAN_CFG4 = 'd0;
localparam CH1_EYESCAN_CFG5 = 'd0;
localparam CH1_EYESCAN_CFG6 = 'd0;
localparam CH1_EYESCAN_CFG7 = 'd0;
localparam CH1_EYESCAN_CFG8 = 'd0;
localparam CH1_EYESCAN_CFG9 = 'd0;
localparam CH1_FABRIC_INTF_CFG0 = 'd4273993723;
localparam CH1_FABRIC_INTF_CFG1 = 'd197632;
localparam CH1_FABRIC_INTF_CFG2 = 'd537919472;
localparam CH1_FABRIC_INTF_CFG3 = 'd786432;
localparam CH1_FABRIC_INTF_CFG4 = 'd20480;
localparam CH1_FABRIC_INTF_CFG5 = 'd25602;
localparam CH1_INSTANTIATED = 'd0;
localparam CH1_MONITOR_CFG = 'd0;
localparam CH1_PIPE_CTRL_CFG0 = 'd262240;
localparam CH1_PIPE_CTRL_CFG1 = 'd2097811;
localparam CH1_PIPE_CTRL_CFG10 = 'd85983215;
localparam CH1_PIPE_CTRL_CFG2 = 'd9950092;
localparam CH1_PIPE_CTRL_CFG3 = 'd1573167;
localparam CH1_PIPE_CTRL_CFG4 = 'd1078198272;
localparam CH1_PIPE_CTRL_CFG5 = 'd2684354560;
localparam CH1_PIPE_CTRL_CFG6 = 'd1007681636;
localparam CH1_PIPE_CTRL_CFG7 = 'd67149834;
localparam CH1_PIPE_CTRL_CFG8 = 'd33554432;
localparam CH1_PIPE_CTRL_CFG9 = 'd0;
localparam CH1_PIPE_TX_EQ_CFG0 = 'd175467487;
localparam CH1_PIPE_TX_EQ_CFG1 = 'd152233553;
localparam CH1_PIPE_TX_EQ_CFG2 = 'd8258;
localparam CH1_PIPE_TX_EQ_CFG3 = 'd393618;
localparam CH1_RESET_BYP_HDSHK_CFG = 'd0;
localparam CH1_RESET_CFG = 'd135266341;
localparam CH1_RESET_LOOPER_ID_CFG = 'd2113632;
localparam CH1_RESET_LOOP_ID_CFG0 = 'd528;
localparam CH1_RESET_LOOP_ID_CFG1 = 'd106181136;
localparam CH1_RESET_LOOP_ID_CFG2 = 'd17185;
localparam CH1_RESET_TIME_CFG0 = 'd34636801;
localparam CH1_RESET_TIME_CFG1 = 'd34636833;
localparam CH1_RESET_TIME_CFG2 = 'd34636833;
localparam CH1_RESET_TIME_CFG3 = 'd2231903265;
localparam CH1_RXOUTCLK_FREQ = 390.625;
localparam CH1_RXOUTCLK_REF_FREQ = 125;
localparam CH1_RXOUTCLK_REF_SOURCE = "HSCLK0_LCPLLGTREFCLK0";
localparam CH1_RX_CDR_CFG0 = 'd3019898946;
localparam CH1_RX_CDR_CFG1 = 'd1610612992;
localparam CH1_RX_CDR_CFG2 = 'd134236777;
localparam CH1_RX_CDR_CFG3 = 'd744694;
localparam CH1_RX_CDR_CFG4 = 'd607924224;
localparam CH1_RX_CRC_CFG0 = 'd30848;
localparam CH1_RX_CRC_CFG1 = 'd505290270;
localparam CH1_RX_CRC_CFG2 = 'd505290270;
localparam CH1_RX_CRC_CFG3 = 'd4294967295;
localparam CH1_RX_CTLE_CFG0 = 'd31195392;
localparam CH1_RX_CTLE_CFG1 = 'd1073741824;
localparam CH1_RX_DACI2V_CFG0 = 'd67145418;
localparam CH1_RX_DFE_CFG0 = 'd3489813512;
localparam CH1_RX_ELASTIC_BUF_CFG0 = 'd2155632704;
localparam CH1_RX_ELASTIC_BUF_CFG1 = 'd2;
localparam CH1_RX_ELASTIC_BUF_CFG2 = 'd0;
localparam CH1_RX_ELASTIC_BUF_CFG3 = 'd2682257408;
localparam CH1_RX_ELASTIC_BUF_CFG4 = 'd0;
localparam CH1_RX_ELASTIC_BUF_CFG5 = 'd0;
localparam CH1_RX_ELASTIC_BUF_CFG6 = 'd4293918720;
localparam CH1_RX_ELASTIC_BUF_CFG7 = 'd67108869;
localparam CH1_RX_ELASTIC_BUF_CFG8 = 'd2033040;
localparam CH1_RX_ELASTIC_BUF_CFG9 = 'd2033040;
localparam CH1_RX_MISC_CFG0 = 'd1342177280;
localparam CH1_RX_OOB_CFG0 = 'd609534468;
localparam CH1_RX_OOB_CFG1 = 'd16925124;
localparam CH1_RX_PAD_CFG0 = 'd0;
localparam CH1_RX_PAD_CFG1 = 'd272910714;
localparam CH1_RX_PCS_CFG0 = 'd674623792;
localparam CH1_RX_PCS_CFG1 = 'd1812204543;
localparam CH1_RX_PCS_CFG2 = 'd1073742049;
localparam CH1_RX_PCS_CFG3 = 'd471666447;
localparam CH1_RX_PCS_CFG4 = 'd1115725826;
localparam CH1_RX_PHALIGN_CFG0 = 'd3;
localparam CH1_RX_PHALIGN_CFG1 = 'd8617984;
localparam CH1_RX_PHALIGN_CFG2 = 'd117248;
localparam CH1_RX_PHALIGN_CFG3 = 'd229376;
localparam CH1_RX_PHALIGN_CFG4 = 'd522;
localparam CH1_RX_PHALIGN_CFG5 = 'd50462720;
localparam CH1_TXOUTCLK_FREQ = 390.625;
localparam CH1_TXOUTCLK_REF_FREQ = 125;
localparam CH1_TXOUTCLK_REF_SOURCE = "HSCLK0_LCPLLGTREFCLK0";
localparam CH1_TX_10G_CFG0 = 'd0;
localparam CH1_TX_10G_CFG1 = 'd1073741824;
localparam CH1_TX_10G_CFG2 = 'd0;
localparam CH1_TX_10G_CFG3 = 'd0;
localparam CH1_TX_ANA_CFG0 = 'd208;
localparam CH1_TX_CRC_CFG0 = 'd30720;
localparam CH1_TX_CRC_CFG1 = 'd505290270;
localparam CH1_TX_CRC_CFG2 = 'd505290270;
localparam CH1_TX_CRC_CFG3 = 'd4294967295;
localparam CH1_TX_DRV_CFG0 = 'd4194304;
localparam CH1_TX_DRV_CFG1 = 'd6144;
localparam CH1_TX_PCS_CFG0 = 'd2187329825;
localparam CH1_TX_PCS_CFG1 = 'd674583932;
localparam CH1_TX_PCS_CFG2 = 'd357954218;
localparam CH1_TX_PCS_CFG3 = 'd1747587;
localparam CH1_TX_PHALIGN_CFG0 = 'd0;
localparam CH1_TX_PHALIGN_CFG1 = 'd290816;
localparam CH1_TX_PHALIGN_CFG2 = 'd229432;
localparam CH1_TX_PHALIGN_CFG3 = 'd0;
localparam CH1_TX_PHALIGN_CFG4 = 'd402653408;
localparam CH1_TX_PHALIGN_CFG5 = 'd128;
localparam CH1_TX_PIPPM_CFG = 'd33554432;
localparam CH1_TX_SER_CFG0 = 'd0;
localparam CH2_ADAPT_APT_CFG = 'd0;
localparam CH2_ADAPT_CAL_CFG = 'd2179884032;
localparam CH2_ADAPT_DFE_CFG = 'd64;
localparam CH2_ADAPT_GC_CFG0 = 'd9441392;
localparam CH2_ADAPT_GC_CFG1 = 'd178259936;
localparam CH2_ADAPT_GC_CFG2 = 'd2097384;
localparam CH2_ADAPT_GC_CFG3 = 'd178258912;
localparam CH2_ADAPT_GEN_CFG0 = 'd1179648;
localparam CH2_ADAPT_GEN_CFG1 = 'd0;
localparam CH2_ADAPT_GEN_CFG2 = 'd2281701375;
localparam CH2_ADAPT_GEN_CFG3 = 'd268435456;
localparam CH2_ADAPT_H01_CFG = 'd18875040;
localparam CH2_ADAPT_H23_CFG = 'd27263392;
localparam CH2_ADAPT_H45_CFG = 'd27263392;
localparam CH2_ADAPT_H67_CFG = 'd27263392;
localparam CH2_ADAPT_H89_CFG = 'd27263392;
localparam CH2_ADAPT_HAB_CFG = 'd27263392;
localparam CH2_ADAPT_HCD_CFG = 'd27263392;
localparam CH2_ADAPT_HEF_CFG = 'd27263904;
localparam CH2_ADAPT_KH_CFG0 = 'd537426239;
localparam CH2_ADAPT_KH_CFG1 = 'd0;
localparam CH2_ADAPT_KH_CFG2 = 'd17312;
localparam CH2_ADAPT_KH_CFG3 = 'd0;
localparam CH2_ADAPT_KH_CFG4 = 'd31648;
localparam CH2_ADAPT_KH_CFG5 = 'd0;
localparam CH2_ADAPT_KL_CFG0 = 'd32928;
localparam CH2_ADAPT_KL_CFG1 = 'd17312;
localparam CH2_ADAPT_LCK_CFG0 = 'd16384;
localparam CH2_ADAPT_LCK_CFG1 = 'd16384;
localparam CH2_ADAPT_LCK_CFG2 = 'd0;
localparam CH2_ADAPT_LCK_CFG3 = 'd0;
localparam CH2_ADAPT_LOP_CFG = 'd3992979040;
localparam CH2_ADAPT_OS_CFG = 'd2147483936;
localparam CH2_CHCLK_ILO_CFG = 'd6553651;
localparam CH2_CHCLK_MISC_CFG = 'd4169260831;
localparam CH2_CHCLK_RSV_CFG = 'd0;
localparam CH2_CHCLK_RXCAL_CFG = 'd138166272;
localparam CH2_CHCLK_RXCAL_CFG1 = 'd0;
localparam CH2_CHCLK_RXCAL_CFG2 = 'd0;
localparam CH2_CHCLK_RXPI_CFG = 'd5244940;
localparam CH2_CHCLK_TXCAL_CFG = 'd4194336;
localparam CH2_CHCLK_TXPI_CFG0 = 'd4655119;
localparam CH2_CHL_RSV_CFG0 = 'd3330277385;
localparam CH2_CHL_RSV_CFG1 = 'd1560;
localparam CH2_CHL_RSV_CFG2 = 'd6227344;
localparam CH2_CHL_RSV_CFG3 = 'd0;
localparam CH2_CHL_RSV_CFG4 = 'd0;
localparam CH2_DA_CFG = 'd655370;
localparam CH2_EYESCAN_CFG0 = 'd2048;
localparam CH2_EYESCAN_CFG1 = 'd0;
localparam CH2_EYESCAN_CFG10 = 'd0;
localparam CH2_EYESCAN_CFG11 = 'd0;
localparam CH2_EYESCAN_CFG12 = 'd0;
localparam CH2_EYESCAN_CFG13 = 'd0;
localparam CH2_EYESCAN_CFG14 = 'd0;
localparam CH2_EYESCAN_CFG15 = 'd0;
localparam CH2_EYESCAN_CFG16 = 'd0;
localparam CH2_EYESCAN_CFG2 = 'd0;
localparam CH2_EYESCAN_CFG3 = 'd0;
localparam CH2_EYESCAN_CFG4 = 'd0;
localparam CH2_EYESCAN_CFG5 = 'd0;
localparam CH2_EYESCAN_CFG6 = 'd0;
localparam CH2_EYESCAN_CFG7 = 'd0;
localparam CH2_EYESCAN_CFG8 = 'd0;
localparam CH2_EYESCAN_CFG9 = 'd0;
localparam CH2_FABRIC_INTF_CFG0 = 'd4273993723;
localparam CH2_FABRIC_INTF_CFG1 = 'd197632;
localparam CH2_FABRIC_INTF_CFG2 = 'd537919472;
localparam CH2_FABRIC_INTF_CFG3 = 'd786432;
localparam CH2_FABRIC_INTF_CFG4 = 'd20480;
localparam CH2_FABRIC_INTF_CFG5 = 'd25602;
localparam CH2_INSTANTIATED = 'd0;
localparam CH2_MONITOR_CFG = 'd0;
localparam CH2_PIPE_CTRL_CFG0 = 'd262240;
localparam CH2_PIPE_CTRL_CFG1 = 'd2097811;
localparam CH2_PIPE_CTRL_CFG10 = 'd85983215;
localparam CH2_PIPE_CTRL_CFG2 = 'd9950092;
localparam CH2_PIPE_CTRL_CFG3 = 'd1573167;
localparam CH2_PIPE_CTRL_CFG4 = 'd1078198272;
localparam CH2_PIPE_CTRL_CFG5 = 'd2684354560;
localparam CH2_PIPE_CTRL_CFG6 = 'd1007681636;
localparam CH2_PIPE_CTRL_CFG7 = 'd67149834;
localparam CH2_PIPE_CTRL_CFG8 = 'd33554432;
localparam CH2_PIPE_CTRL_CFG9 = 'd0;
localparam CH2_PIPE_TX_EQ_CFG0 = 'd175467487;
localparam CH2_PIPE_TX_EQ_CFG1 = 'd152233553;
localparam CH2_PIPE_TX_EQ_CFG2 = 'd8258;
localparam CH2_PIPE_TX_EQ_CFG3 = 'd393618;
localparam CH2_RESET_BYP_HDSHK_CFG = 'd0;
localparam CH2_RESET_CFG = 'd135266341;
localparam CH2_RESET_LOOPER_ID_CFG = 'd2113632;
localparam CH2_RESET_LOOP_ID_CFG0 = 'd528;
localparam CH2_RESET_LOOP_ID_CFG1 = 'd106181136;
localparam CH2_RESET_LOOP_ID_CFG2 = 'd17185;
localparam CH2_RESET_TIME_CFG0 = 'd34636801;
localparam CH2_RESET_TIME_CFG1 = 'd34636833;
localparam CH2_RESET_TIME_CFG2 = 'd34636833;
localparam CH2_RESET_TIME_CFG3 = 'd2231903265;
localparam CH2_RXOUTCLK_FREQ = 390.625;
localparam CH2_RXOUTCLK_REF_FREQ = 100;
localparam CH2_RXOUTCLK_REF_SOURCE = "HSCLK1_LCPLLGTREFCLK0";
localparam CH2_RX_CDR_CFG0 = 'd3019898946;
localparam CH2_RX_CDR_CFG1 = 'd1610612992;
localparam CH2_RX_CDR_CFG2 = 'd134236777;
localparam CH2_RX_CDR_CFG3 = 'd744694;
localparam CH2_RX_CDR_CFG4 = 'd607924224;
localparam CH2_RX_CRC_CFG0 = 'd30848;
localparam CH2_RX_CRC_CFG1 = 'd505290270;
localparam CH2_RX_CRC_CFG2 = 'd505290270;
localparam CH2_RX_CRC_CFG3 = 'd4294967295;
localparam CH2_RX_CTLE_CFG0 = 'd31195392;
localparam CH2_RX_CTLE_CFG1 = 'd1073741824;
localparam CH2_RX_DACI2V_CFG0 = 'd67145418;
localparam CH2_RX_DFE_CFG0 = 'd3489813512;
localparam CH2_RX_ELASTIC_BUF_CFG0 = 'd2155632704;
localparam CH2_RX_ELASTIC_BUF_CFG1 = 'd2;
localparam CH2_RX_ELASTIC_BUF_CFG2 = 'd0;
localparam CH2_RX_ELASTIC_BUF_CFG3 = 'd2682257408;
localparam CH2_RX_ELASTIC_BUF_CFG4 = 'd0;
localparam CH2_RX_ELASTIC_BUF_CFG5 = 'd0;
localparam CH2_RX_ELASTIC_BUF_CFG6 = 'd4293918720;
localparam CH2_RX_ELASTIC_BUF_CFG7 = 'd67108869;
localparam CH2_RX_ELASTIC_BUF_CFG8 = 'd2033040;
localparam CH2_RX_ELASTIC_BUF_CFG9 = 'd2033040;
localparam CH2_RX_MISC_CFG0 = 'd1342177280;
localparam CH2_RX_OOB_CFG0 = 'd609534468;
localparam CH2_RX_OOB_CFG1 = 'd16925124;
localparam CH2_RX_PAD_CFG0 = 'd0;
localparam CH2_RX_PAD_CFG1 = 'd272910714;
localparam CH2_RX_PCS_CFG0 = 'd674623792;
localparam CH2_RX_PCS_CFG1 = 'd1812204543;
localparam CH2_RX_PCS_CFG2 = 'd1073742049;
localparam CH2_RX_PCS_CFG3 = 'd471666447;
localparam CH2_RX_PCS_CFG4 = 'd1115725826;
localparam CH2_RX_PHALIGN_CFG0 = 'd3;
localparam CH2_RX_PHALIGN_CFG1 = 'd8617984;
localparam CH2_RX_PHALIGN_CFG2 = 'd117248;
localparam CH2_RX_PHALIGN_CFG3 = 'd229376;
localparam CH2_RX_PHALIGN_CFG4 = 'd522;
localparam CH2_RX_PHALIGN_CFG5 = 'd50462720;
localparam CH2_TXOUTCLK_FREQ = 390.625;
localparam CH2_TXOUTCLK_REF_FREQ = 100;
localparam CH2_TXOUTCLK_REF_SOURCE = "HSCLK1_LCPLLGTREFCLK0";
localparam CH2_TX_10G_CFG0 = 'd0;
localparam CH2_TX_10G_CFG1 = 'd1073741824;
localparam CH2_TX_10G_CFG2 = 'd0;
localparam CH2_TX_10G_CFG3 = 'd0;
localparam CH2_TX_ANA_CFG0 = 'd208;
localparam CH2_TX_CRC_CFG0 = 'd30720;
localparam CH2_TX_CRC_CFG1 = 'd505290270;
localparam CH2_TX_CRC_CFG2 = 'd505290270;
localparam CH2_TX_CRC_CFG3 = 'd4294967295;
localparam CH2_TX_DRV_CFG0 = 'd4194304;
localparam CH2_TX_DRV_CFG1 = 'd6144;
localparam CH2_TX_PCS_CFG0 = 'd2187329825;
localparam CH2_TX_PCS_CFG1 = 'd674583932;
localparam CH2_TX_PCS_CFG2 = 'd357954218;
localparam CH2_TX_PCS_CFG3 = 'd1747587;
localparam CH2_TX_PHALIGN_CFG0 = 'd0;
localparam CH2_TX_PHALIGN_CFG1 = 'd290816;
localparam CH2_TX_PHALIGN_CFG2 = 'd229432;
localparam CH2_TX_PHALIGN_CFG3 = 'd0;
localparam CH2_TX_PHALIGN_CFG4 = 'd402653408;
localparam CH2_TX_PHALIGN_CFG5 = 'd128;
localparam CH2_TX_PIPPM_CFG = 'd33554432;
localparam CH2_TX_SER_CFG0 = 'd0;
localparam CH3_ADAPT_APT_CFG = 'd0;
localparam CH3_ADAPT_CAL_CFG = 'd2179884032;
localparam CH3_ADAPT_DFE_CFG = 'd64;
localparam CH3_ADAPT_GC_CFG0 = 'd9441392;
localparam CH3_ADAPT_GC_CFG1 = 'd178259936;
localparam CH3_ADAPT_GC_CFG2 = 'd2097384;
localparam CH3_ADAPT_GC_CFG3 = 'd178258912;
localparam CH3_ADAPT_GEN_CFG0 = 'd1179648;
localparam CH3_ADAPT_GEN_CFG1 = 'd0;
localparam CH3_ADAPT_GEN_CFG2 = 'd2281701375;
localparam CH3_ADAPT_GEN_CFG3 = 'd268435456;
localparam CH3_ADAPT_H01_CFG = 'd18875040;
localparam CH3_ADAPT_H23_CFG = 'd27263392;
localparam CH3_ADAPT_H45_CFG = 'd27263392;
localparam CH3_ADAPT_H67_CFG = 'd27263392;
localparam CH3_ADAPT_H89_CFG = 'd27263392;
localparam CH3_ADAPT_HAB_CFG = 'd27263392;
localparam CH3_ADAPT_HCD_CFG = 'd27263392;
localparam CH3_ADAPT_HEF_CFG = 'd27263904;
localparam CH3_ADAPT_KH_CFG0 = 'd537426239;
localparam CH3_ADAPT_KH_CFG1 = 'd0;
localparam CH3_ADAPT_KH_CFG2 = 'd17312;
localparam CH3_ADAPT_KH_CFG3 = 'd0;
localparam CH3_ADAPT_KH_CFG4 = 'd31648;
localparam CH3_ADAPT_KH_CFG5 = 'd0;
localparam CH3_ADAPT_KL_CFG0 = 'd32928;
localparam CH3_ADAPT_KL_CFG1 = 'd17312;
localparam CH3_ADAPT_LCK_CFG0 = 'd16384;
localparam CH3_ADAPT_LCK_CFG1 = 'd16384;
localparam CH3_ADAPT_LCK_CFG2 = 'd0;
localparam CH3_ADAPT_LCK_CFG3 = 'd0;
localparam CH3_ADAPT_LOP_CFG = 'd3992979040;
localparam CH3_ADAPT_OS_CFG = 'd2147483936;
localparam CH3_CHCLK_ILO_CFG = 'd6553651;
localparam CH3_CHCLK_MISC_CFG = 'd4169260831;
localparam CH3_CHCLK_RSV_CFG = 'd0;
localparam CH3_CHCLK_RXCAL_CFG = 'd138166272;
localparam CH3_CHCLK_RXCAL_CFG1 = 'd0;
localparam CH3_CHCLK_RXCAL_CFG2 = 'd0;
localparam CH3_CHCLK_RXPI_CFG = 'd5244940;
localparam CH3_CHCLK_TXCAL_CFG = 'd4194336;
localparam CH3_CHCLK_TXPI_CFG0 = 'd4655119;
localparam CH3_CHL_RSV_CFG0 = 'd3330277385;
localparam CH3_CHL_RSV_CFG1 = 'd1560;
localparam CH3_CHL_RSV_CFG2 = 'd6227344;
localparam CH3_CHL_RSV_CFG3 = 'd0;
localparam CH3_CHL_RSV_CFG4 = 'd0;
localparam CH3_DA_CFG = 'd655370;
localparam CH3_EYESCAN_CFG0 = 'd2048;
localparam CH3_EYESCAN_CFG1 = 'd0;
localparam CH3_EYESCAN_CFG10 = 'd0;
localparam CH3_EYESCAN_CFG11 = 'd0;
localparam CH3_EYESCAN_CFG12 = 'd0;
localparam CH3_EYESCAN_CFG13 = 'd0;
localparam CH3_EYESCAN_CFG14 = 'd0;
localparam CH3_EYESCAN_CFG15 = 'd0;
localparam CH3_EYESCAN_CFG16 = 'd0;
localparam CH3_EYESCAN_CFG2 = 'd0;
localparam CH3_EYESCAN_CFG3 = 'd0;
localparam CH3_EYESCAN_CFG4 = 'd0;
localparam CH3_EYESCAN_CFG5 = 'd0;
localparam CH3_EYESCAN_CFG6 = 'd0;
localparam CH3_EYESCAN_CFG7 = 'd0;
localparam CH3_EYESCAN_CFG8 = 'd0;
localparam CH3_EYESCAN_CFG9 = 'd0;
localparam CH3_FABRIC_INTF_CFG0 = 'd4273993723;
localparam CH3_FABRIC_INTF_CFG1 = 'd1024;
localparam CH3_FABRIC_INTF_CFG2 = 'd537919472;
localparam CH3_FABRIC_INTF_CFG3 = 'd0;
localparam CH3_FABRIC_INTF_CFG4 = 'd20480;
localparam CH3_FABRIC_INTF_CFG5 = 'd25602;
localparam CH3_INSTANTIATED = 'd1;
localparam CH3_MONITOR_CFG = 'd0;
localparam CH3_PIPE_CTRL_CFG0 = 'd262240;
localparam CH3_PIPE_CTRL_CFG1 = 'd2097811;
localparam CH3_PIPE_CTRL_CFG10 = 'd85983215;
localparam CH3_PIPE_CTRL_CFG2 = 'd9950092;
localparam CH3_PIPE_CTRL_CFG3 = 'd77070639;
localparam CH3_PIPE_CTRL_CFG4 = 'd4456448;
localparam CH3_PIPE_CTRL_CFG5 = 'd2684354560;
localparam CH3_PIPE_CTRL_CFG6 = 'd1007681636;
localparam CH3_PIPE_CTRL_CFG7 = 'd67149834;
localparam CH3_PIPE_CTRL_CFG8 = 'd33677432;
localparam CH3_PIPE_CTRL_CFG9 = 'd0;
localparam CH3_PIPE_TX_EQ_CFG0 = 'd175467487;
localparam CH3_PIPE_TX_EQ_CFG1 = 'd152233553;
localparam CH3_PIPE_TX_EQ_CFG2 = 'd8258;
localparam CH3_PIPE_TX_EQ_CFG3 = 'd393618;
localparam CH3_RESET_BYP_HDSHK_CFG = 'd0;
localparam CH3_RESET_CFG = 'd135266357;
localparam CH3_RESET_LOOPER_ID_CFG = 'd2113632;
localparam CH3_RESET_LOOP_ID_CFG0 = 'd528;
localparam CH3_RESET_LOOP_ID_CFG1 = 'd106181136;
localparam CH3_RESET_LOOP_ID_CFG2 = 'd17185;
localparam CH3_RESET_TIME_CFG0 = 'd34636801;
localparam CH3_RESET_TIME_CFG1 = 'd34636833;
localparam CH3_RESET_TIME_CFG2 = 'd34636833;
localparam CH3_RESET_TIME_CFG3 = 'd2231903265;
localparam CH3_RXOUTCLK_FREQ = 150;
localparam CH3_RXOUTCLK_REF_FREQ = 100;
localparam CH3_RXOUTCLK_REF_SOURCE = "HSCLK1_LCPLLGTREFCLK0";
localparam CH3_RX_CDR_CFG0 = 'd2885681218;
localparam CH3_RX_CDR_CFG1 = 'd1610612992;
localparam CH3_RX_CDR_CFG2 = 'd134236745;
localparam CH3_RX_CDR_CFG3 = 'd744694;
localparam CH3_RX_CDR_CFG4 = 'd607924224;
localparam CH3_RX_CRC_CFG0 = 'd30848;
localparam CH3_RX_CRC_CFG1 = 'd505290270;
localparam CH3_RX_CRC_CFG2 = 'd505290270;
localparam CH3_RX_CRC_CFG3 = 'd4294967295;
localparam CH3_RX_CTLE_CFG0 = 'd31195392;
localparam CH3_RX_CTLE_CFG1 = 'd1073741824;
localparam CH3_RX_DACI2V_CFG0 = 'd67145418;
localparam CH3_RX_DFE_CFG0 = 'd3489813512;
localparam CH3_RX_ELASTIC_BUF_CFG0 = 'd4202594;
localparam CH3_RX_ELASTIC_BUF_CFG1 = 'd533522418;
localparam CH3_RX_ELASTIC_BUF_CFG2 = 'd3221225599;
localparam CH3_RX_ELASTIC_BUF_CFG3 = 'd3755999232;
localparam CH3_RX_ELASTIC_BUF_CFG4 = 'd0;
localparam CH3_RX_ELASTIC_BUF_CFG5 = 'd0;
localparam CH3_RX_ELASTIC_BUF_CFG6 = 'd4293918720;
localparam CH3_RX_ELASTIC_BUF_CFG7 = 'd67108868;
localparam CH3_RX_ELASTIC_BUF_CFG8 = 'd2033040;
localparam CH3_RX_ELASTIC_BUF_CFG9 = 'd2033040;
localparam CH3_RX_MISC_CFG0 = 'd1342177281;
localparam CH3_RX_OOB_CFG0 = 'd609534468;
localparam CH3_RX_OOB_CFG1 = 'd16925124;
localparam CH3_RX_PAD_CFG0 = 'd0;
localparam CH3_RX_PAD_CFG1 = 'd272910714;
localparam CH3_RX_PCS_CFG0 = 'd3895849135;
localparam CH3_RX_PCS_CFG1 = 'd605036671;
localparam CH3_RX_PCS_CFG2 = 'd1074118912;
localparam CH3_RX_PCS_CFG3 = 'd471666447;
localparam CH3_RX_PCS_CFG4 = 'd3263209474;
localparam CH3_RX_PHALIGN_CFG0 = 'd3;
localparam CH3_RX_PHALIGN_CFG1 = 'd8617984;
localparam CH3_RX_PHALIGN_CFG2 = 'd117248;
localparam CH3_RX_PHALIGN_CFG3 = 'd229376;
localparam CH3_RX_PHALIGN_CFG4 = 'd522;
localparam CH3_RX_PHALIGN_CFG5 = 'd50462720;
localparam CH3_TXOUTCLK_FREQ = 150;
localparam CH3_TXOUTCLK_REF_FREQ = 100;
localparam CH3_TXOUTCLK_REF_SOURCE = "HSCLK1_LCPLLGTREFCLK0";
localparam CH3_TX_10G_CFG0 = 'd0;
localparam CH3_TX_10G_CFG1 = 'd1073741824;
localparam CH3_TX_10G_CFG2 = 'd0;
localparam CH3_TX_10G_CFG3 = 'd0;
localparam CH3_TX_ANA_CFG0 = 'd208;
localparam CH3_TX_CRC_CFG0 = 'd30720;
localparam CH3_TX_CRC_CFG1 = 'd505290270;
localparam CH3_TX_CRC_CFG2 = 'd505290270;
localparam CH3_TX_CRC_CFG3 = 'd4294967295;
localparam CH3_TX_DRV_CFG0 = 'd4194304;
localparam CH3_TX_DRV_CFG1 = 'd6144;
localparam CH3_TX_PCS_CFG0 = 'd559022336;
localparam CH3_TX_PCS_CFG1 = 'd674583932;
localparam CH3_TX_PCS_CFG2 = 'd357954218;
localparam CH3_TX_PCS_CFG3 = 'd1747587;
localparam CH3_TX_PHALIGN_CFG0 = 'd0;
localparam CH3_TX_PHALIGN_CFG1 = 'd290816;
localparam CH3_TX_PHALIGN_CFG2 = 'd229432;
localparam CH3_TX_PHALIGN_CFG3 = 'd0;
localparam CH3_TX_PHALIGN_CFG4 = 'd402653408;
localparam CH3_TX_PHALIGN_CFG5 = 'd160;
localparam CH3_TX_PIPPM_CFG = 'd33554432;
localparam CH3_TX_SER_CFG0 = 'd0;
localparam CTRL_RSV_CFG0 = 'd30744;
localparam CTRL_RSV_CFG1 = 'd0;
localparam HS0_LCPLL_IPS_PIN_EN = 'd0;
localparam HS0_LCPLL_IPS_REFCLK_SEL = 'd1;
localparam HS0_LCPLL_REFCLK_MAP0  = 'd0;
localparam HS0_LCPLL_REFCLK_MAP1  = 'd1;
localparam HS0_LCPLL_REFCLK_MAP2  = 'd2;
localparam HS0_LCPLL_REFCLK_MAP3  = 'd3;
localparam HS0_LCPLL_REFCLK_MAP4  = 'd4;
localparam HS0_LCPLL_REFCLK_MAP5  = 'd5;
localparam HS0_LCPLL_REFCLK_MAP6  = 'd6;
localparam HS0_LCPLL_REFCLK_MAP7  = 'd7;
localparam HS0_RPLL_IPS_PIN_EN = 'd0;
localparam HS0_RPLL_IPS_REFCLK_SEL = 'd1;
localparam HS0_RPLL_REFCLK_MAP0  = 'd0;
localparam HS0_RPLL_REFCLK_MAP1  = 'd1;
localparam HS0_RPLL_REFCLK_MAP2  = 'd2;
localparam HS0_RPLL_REFCLK_MAP3  = 'd3;
localparam HS0_RPLL_REFCLK_MAP4  = 'd4;
localparam HS0_RPLL_REFCLK_MAP5  = 'd5;
localparam HS0_RPLL_REFCLK_MAP6  = 'd6;
localparam HS0_RPLL_REFCLK_MAP7  = 'd7;
localparam HS1_LCPLL_IPS_PIN_EN = 'd0;
localparam HS1_LCPLL_IPS_REFCLK_SEL = 'd1;
localparam HS1_LCPLL_REFCLK_MAP0  = 'd0;
localparam HS1_LCPLL_REFCLK_MAP1  = 'd2;
localparam HS1_LCPLL_REFCLK_MAP2  = 'd1;
localparam HS1_LCPLL_REFCLK_MAP3  = 'd3;
localparam HS1_LCPLL_REFCLK_MAP4  = 'd4;
localparam HS1_LCPLL_REFCLK_MAP5  = 'd5;
localparam HS1_LCPLL_REFCLK_MAP6  = 'd6;
localparam HS1_LCPLL_REFCLK_MAP7  = 'd7;
localparam HS1_RPLL_IPS_PIN_EN = 'd0;
localparam HS1_RPLL_IPS_REFCLK_SEL = 'd1;
localparam HS1_RPLL_REFCLK_MAP0  = 'd0;
localparam HS1_RPLL_REFCLK_MAP1  = 'd2;
localparam HS1_RPLL_REFCLK_MAP2  = 'd1;
localparam HS1_RPLL_REFCLK_MAP3  = 'd3;
localparam HS1_RPLL_REFCLK_MAP4  = 'd4;
localparam HS1_RPLL_REFCLK_MAP5  = 'd5;
localparam HS1_RPLL_REFCLK_MAP6  = 'd6;
localparam HS1_RPLL_REFCLK_MAP7  = 'd7;
localparam HSCLK0_HSDIST_CFG = 'd30;
localparam HSCLK0_INSTANTIATED = 'd0;
localparam HSCLK0_LCPLL_CFG0 = 'd4210436;
localparam HSCLK0_LCPLL_CFG1 = 'd68701952;
localparam HSCLK0_LCPLL_CFG2 = 'd2185429512;
localparam HSCLK0_LCPLL_LGC_CFG0 = 'd3855911696;
localparam HSCLK0_LCPLL_LGC_CFG1 = 'd2484213888;
localparam HSCLK0_LCPLL_LGC_CFG2 = 'd1114385;
localparam HSCLK0_RPLL_CFG0 = 'd2147516356;
localparam HSCLK0_RPLL_CFG1 = 'd132267816;
localparam HSCLK0_RPLL_CFG2 = 'd11740105;
localparam HSCLK0_RPLL_LGC_CFG0 = 'd3855912336;
localparam HSCLK0_RPLL_LGC_CFG1 = 'd2484213888;
localparam HSCLK0_RPLL_LGC_CFG2 = 'd1114385;
localparam HSCLK1_HSDIST_CFG = 'd65566;
localparam HSCLK1_INSTANTIATED = 'd1;
localparam HSCLK1_LCPLL_CFG0 = 'd4210436;
localparam HSCLK1_LCPLL_CFG1 = 'd68701952;
localparam HSCLK1_LCPLL_CFG2 = 'd2184970760;
localparam HSCLK1_LCPLL_LGC_CFG0 = 'd3855911696;
localparam HSCLK1_LCPLL_LGC_CFG1 = 'd2484213888;
localparam HSCLK1_LCPLL_LGC_CFG2 = 'd1114385;
localparam HSCLK1_RPLL_CFG0 = 'd2147516356;
localparam HSCLK1_RPLL_CFG1 = 'd132267816;
localparam HSCLK1_RPLL_CFG2 = 'd11740105;
localparam HSCLK1_RPLL_LGC_CFG0 = 'd3855912336;
localparam HSCLK1_RPLL_LGC_CFG1 = 'd2484213888;
localparam HSCLK1_RPLL_LGC_CFG2 = 'd1114385;
localparam MST_RESET_CFG = 'd2320667656;
localparam PIN_CFG0 = 'd8929817;
localparam POR_CFG = 'd285440;
localparam QUAD_INSTANTIATED = 'd1;
localparam RCALBG0_CFG0 = 'd976;
localparam RCALBG0_CFG1 = 'd64;
localparam RCALBG0_CFG2 = 'd0;
localparam RCALBG0_CFG3 = 'd2147483650;
localparam RCALBG0_CFG4 = 'd279;
localparam RCALBG0_CFG5 = 'd691;
localparam RCALBG1_CFG0 = 'd976;
localparam RCALBG1_CFG1 = 'd64;
localparam RCALBG1_CFG2 = 'd0;
localparam RCALBG1_CFG3 = 'd2147483650;
localparam RCALBG1_CFG4 = 'd279;
localparam RCALBG1_CFG5 = 'd691;
localparam RXRSTDONE_DIST_SEL = 'd0;
localparam STAT_NPI_REG_LIST = "3000:3004,3010:3014,3020:3024,3034:304C,3070:3098,30A8:30B4,30BC:30EC,30F4:3178,3180:3184,318C:3190,3198:31A0,31B0:31D8,31E0:31E8,31F0:3228,3230:3264,326C:3274,3280,3294:329C,32A8,32BC:32E4,32FC,3430:3444,344C,3470:3498,34A8:34B4,34BC:34EC,34F4:3578,3580:3584,358C:3590,3598:35A0,35B0:35D8,35E0:35E8,35F0:3628,3630:3664,366C:3674,3680,3694:369C,36A8,36BC:36E4,3834:383C,3848,3870:3898,38A8:38B4,38BC:38EC,38F4:3978,3980:3984,398C:3990,3998:39A0,39B0:39D8,39E0:39E8,39F0:3A28,3A30:3A64,3A6C:3A74,3A80,3A94:3A9C,3AA8,3ABC:3AE4,3AFC,3C08,3C30:3C3C,3C48:3C4C,3C70:3C98,3CA8:3CB4,3CBC:3CEC,3CF4:3D78,3D80:3D84,3D8C:3D90,3D98:3DA0,3DB0:3DD8,3DE0:3DE8,3DF0:3E28,3E30:3E64,3E6C:3E74,3E80,3E94:3E9C,3EA8,3EBC:3EE4";
localparam TERMPROG_CFG = 'd0;
localparam TXRSTDONE_DIST_SEL = 'd0;
localparam UB_CFG0 = 'd1933574144;
localparam CH0_SIM_MODE = "FAST";
localparam CH0_SIM_RECEIVER_DETECT_PASS = "TRUE";
localparam CH0_SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
localparam CH1_SIM_MODE = "FAST";
localparam CH1_SIM_RECEIVER_DETECT_PASS = "TRUE";
localparam CH1_SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
localparam CH2_SIM_MODE = "FAST";
localparam CH2_SIM_RECEIVER_DETECT_PASS = "TRUE";
localparam CH2_SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
localparam CH3_SIM_MODE = "FAST";
localparam CH3_SIM_RECEIVER_DETECT_PASS = "TRUE";
localparam CH3_SIM_TX_EIDLE_DRIVE_LEVEL = "Z";
localparam QUAD_SIM_MODE = "FAST";
localparam QUAD_SIM_RESET_SPEEDUP = "TRUE";
localparam CH3_SIM_RESET_SPEEDUP = "TRUE";
localparam CH2_SIM_RESET_SPEEDUP = "TRUE";
localparam CH1_SIM_RESET_SPEEDUP = "TRUE";
localparam CH0_SIM_RESET_SPEEDUP = "TRUE";
localparam SIM_DEVICE = "";
localparam MEMORY_INIT_FILE = "extended_phy_layer_gtwiz_versal_0_0_gt_quad_base_0.mem";
localparam SIM_VERSION = "2";
