// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_BFR_MATMULX_DEFINES_VH
`else
`define B_BFR_MATMULX_DEFINES_VH

// Look-up table parameters
//

`define BFR_MATMULX_ADDR_N  7
`define BFR_MATMULX_ADDR_SZ 32
`define BFR_MATMULX_DATA_SZ 64

// Attribute addresses
//

`define BFR_MATMULX__ACTIVE_DUTYCYCLE    32'h00000000
`define BFR_MATMULX__ACTIVE_DUTYCYCLE_SZ 64

`define BFR_MATMULX__BFRTYPE    32'h00000001
`define BFR_MATMULX__BFRTYPE_SZ 56

`define BFR_MATMULX__CLK_FREQ    32'h00000002
`define BFR_MATMULX__CLK_FREQ_SZ 64

`define BFR_MATMULX__EN_CLK_DOUBLER    32'h00000003
`define BFR_MATMULX__EN_CLK_DOUBLER_SZ 1

`define BFR_MATMULX__NUM_COMPUTE    32'h00000004
`define BFR_MATMULX__NUM_COMPUTE_SZ 4

`define BFR_MATMULX__NUM_MEMORY    32'h00000005
`define BFR_MATMULX__NUM_MEMORY_SZ 4

`define BFR_MATMULX__XPA_CFG0    32'h00000006
`define BFR_MATMULX__XPA_CFG0_SZ 16

`endif  // B_BFR_MATMULX_DEFINES_VH