----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module checks the validity of the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_desencapsulation is
  generic (
    G_VC_NUM       : integer := 8                                                  --! Number of virtual channel
 );
  port (
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- DBUFI interface
    RD_DATA_DBUFI          : in std_logic_vector(36-1 downto 0);    -- Data read bus
    RD_DATA_EN_DBUFI       : out  std_logic;                                -- Read command
    RD_DATA_VLD_DBUFI      : in std_logic;                                -- Data valid
    -- DOBUF interface
    FCT_FAR_END_DDES       : out  std_logic_vector(G_VC_NUM-1 downto 0);    -- Data write bus
    WR_MULT                : out  vc_multiplier(G_VC_NUM-1 downto 0);
    -- DIBUF interface
    WR_DATA_DDES           : out  vc_data_k_array(G_VC_NUM downto 0);    -- Data write vc & broadcast
    WR_DATA_EN_DDES        : out  std_logic_vector(G_VC_NUM downto 0)   -- Write command vc & broadcast
  );
end data_desencapsulation;

architecture rtl of data_desencapsulation is
---------------------------------------------------------
-----                  Declaration signals          -----
---------------------------------------------------------
constant C_DATA_DBUFI_WIDTH : integer := 36; -- a mettre dans pkg
constant C_BYTE_WIDTH : integer := 8;
-- valeur a changer
constant C_D16_2_SYMB : std_logic_vector(07 downto 00) := x"FA";  --! D16.2 SDF
constant C_D29_2_SYMB : std_logic_vector(07 downto 00) := x"FB";  --! D29.2 SBF

signal data_detected      : std_logic; --high when sdf read
signal broadcast_detected : std_logic; --high when sbf read
signal vc_nb              : integer;    

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_desencapsulation
-- Description: desencapsulate each frame 
---------------------------------------------------------
p_desencapsulation : process(CLK, RST_N)     
begin
  if RST_N = '0' then
    FCT_FAR_END_DDES           <= (others => '0'); 
    WR_DATA_DDES               <= (others =>(others => '0'));
    WR_MULT                    <= (others =>(others => '0'));
    WR_DATA_EN_DDES            <= (others => '0');
    RD_DATA_EN_DBUFI           <= '0';
    data_detected              <= '0';
    broadcast_detected         <= '0';
  elsif rising_edge(CLK) then
    RD_DATA_EN_DBUFI       <= '1';
    if RD_DATA_VLD_DBUFI = '1' then
      --                      msb = 35
      if RD_DATA_DBUFI(C_DATA_DBUFI_WIDTH - 3 downto C_DATA_DBUFI_WIDTH - 4) = "01" then --reading a K character
        --                              15 downto 0
        if RD_DATA_DBUFI(C_BYTE_WIDTH*2 - 1 downto 0) =  C_D16_2_SYMB & C_K28_7_SYMB  then -- SDF
          data_detected                                 <= '1';
          vc_nb                                         <= to_integer(unsigned(RD_DATA_DBUFI(C_BYTE_WIDTH*3 -1 downto C_BYTE_WIDTH*2)));
        --                                 15 downto 0
        elsif RD_DATA_DBUFI(C_BYTE_WIDTH*2 - 1 downto 0) =  C_D29_2_SYMB & C_K28_7_SYMB then --SBF
          broadcast_detected                            <= '1';
        --                                 7 downto 0
        elsif RD_DATA_DBUFI(C_BYTE_WIDTH - 1 downto 0) = C_K28_3_SYMB then --FCT
          --                                                       12 downto 8                                                          23 downto 21
          WR_MULT(to_integer(unsigned(RD_DATA_DBUFI(C_BYTE_WIDTH +4 downto C_BYTE_WIDTH)))) <= std_logic_vector(to_unsigned(to_integer(unsigned(RD_DATA_DBUFI(C_BYTE_WIDTH*2 -1 downto C_BYTE_WIDTH*2 - 3)))+1,4));
          FCT_FAR_END_DDES (to_integer(unsigned(RD_DATA_DBUFI(C_BYTE_WIDTH*2 +4 downto C_BYTE_WIDTH*2)))) <= '1';

        elsif RD_DATA_DBUFI(C_BYTE_WIDTH - 1 downto 0) = C_K28_0_SYMB then --EDF
          data_detected                                 <= '0';
          WR_DATA_EN_DDES                               <= (others => '0');
        elsif RD_DATA_DBUFI(C_BYTE_WIDTH - 1 downto 0) = C_K28_2_SYMB then --EBF
          broadcast_detected                            <= '0';
          WR_DATA_EN_DDES                               <= (others => '0');
        end if;
      else --just normal data
        if data_detected = '1' or broadcast_detected = '1' then 
          if broadcast_detected = '1' then
            WR_DATA_DDES   (G_VC_NUM) <= RD_DATA_DBUFI(C_DATA_DBUFI_WIDTH-1 downto 0);
            WR_DATA_EN_DDES(G_VC_NUM) <= '1';
          else
            WR_DATA_DDES   (vc_nb)      <= RD_DATA_DBUFI(C_DATA_DBUFI_WIDTH-1 downto 0);
            WR_DATA_EN_DDES(vc_nb)      <= '1';
          end if;
        end if;
      end if;
    else --not valid 
      FCT_FAR_END_DDES           <= (others => '0'); 
      WR_DATA_DDES               <= (others =>(others => '0'));
      WR_MULT                    <= (others =>(others => '0'));
      WR_DATA_EN_DDES            <= (others => '0');
    end if;
  end if;
end process;

end architecture rtl;