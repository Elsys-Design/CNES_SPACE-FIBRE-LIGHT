// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_XRAM_DEFINES_VH
`else
`define B_XRAM_DEFINES_VH

// Look-up table parameters
//

`define XRAM_ADDR_N  19
`define XRAM_ADDR_SZ 32
`define XRAM_DATA_SZ 64

// Attribute addresses
//

`define XRAM__MEM_FREQ    32'h00000000
`define XRAM__MEM_FREQ_SZ 64

`define XRAM__PL_INTERFACE_1_FREQUENCY    32'h00000001
`define XRAM__PL_INTERFACE_1_FREQUENCY_SZ 64

`define XRAM__PL_INTERFACE_1_INTERFACE_BANDWIDTH    32'h00000002
`define XRAM__PL_INTERFACE_1_INTERFACE_BANDWIDTH_SZ 15

`define XRAM__PL_INTERFACE_1_INTERFACE_USAGE    32'h00000003
`define XRAM__PL_INTERFACE_1_INTERFACE_USAGE_SZ 1

`define XRAM__PL_INTERFACE_1_INTERFACE_WIDTH    32'h00000004
`define XRAM__PL_INTERFACE_1_INTERFACE_WIDTH_SZ 9

`define XRAM__PL_INTERFACE_1_NUM_MEM_BANKS    32'h00000005
`define XRAM__PL_INTERFACE_1_NUM_MEM_BANKS_SZ 3

`define XRAM__PL_INTERFACE_2_FREQUENCY    32'h00000006
`define XRAM__PL_INTERFACE_2_FREQUENCY_SZ 64

`define XRAM__PL_INTERFACE_2_INTERFACE_BANDWIDTH    32'h00000007
`define XRAM__PL_INTERFACE_2_INTERFACE_BANDWIDTH_SZ 15

`define XRAM__PL_INTERFACE_2_INTERFACE_USAGE    32'h00000008
`define XRAM__PL_INTERFACE_2_INTERFACE_USAGE_SZ 1

`define XRAM__PL_INTERFACE_2_INTERFACE_WIDTH    32'h00000009
`define XRAM__PL_INTERFACE_2_INTERFACE_WIDTH_SZ 9

`define XRAM__PL_INTERFACE_2_NUM_MEM_BANKS    32'h0000000a
`define XRAM__PL_INTERFACE_2_NUM_MEM_BANKS_SZ 3

`define XRAM__PL_INTERFACE_3_FREQUENCY    32'h0000000b
`define XRAM__PL_INTERFACE_3_FREQUENCY_SZ 64

`define XRAM__PL_INTERFACE_3_INTERFACE_BANDWIDTH    32'h0000000c
`define XRAM__PL_INTERFACE_3_INTERFACE_BANDWIDTH_SZ 15

`define XRAM__PL_INTERFACE_3_INTERFACE_USAGE    32'h0000000d
`define XRAM__PL_INTERFACE_3_INTERFACE_USAGE_SZ 1

`define XRAM__PL_INTERFACE_3_INTERFACE_WIDTH    32'h0000000e
`define XRAM__PL_INTERFACE_3_INTERFACE_WIDTH_SZ 9

`define XRAM__PL_INTERFACE_3_NUM_MEM_BANKS    32'h0000000f
`define XRAM__PL_INTERFACE_3_NUM_MEM_BANKS_SZ 3

`define XRAM__PS_INTERFACE_BANDWIDTH    32'h00000010
`define XRAM__PS_INTERFACE_BANDWIDTH_SZ 15

`define XRAM__PS_INTERFACE_NUM_MEM_BANKS    32'h00000011
`define XRAM__PS_INTERFACE_NUM_MEM_BANKS_SZ 3

`define XRAM__PS_INTERFACE_USAGE    32'h00000012
`define XRAM__PS_INTERFACE_USAGE_SZ 1

`endif  // B_XRAM_DEFINES_VH