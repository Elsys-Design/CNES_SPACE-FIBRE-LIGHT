// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTF_COMMON_DEFINES_VH
`else
`define B_GTF_COMMON_DEFINES_VH

// Look-up table parameters
//

`define GTF_COMMON_ADDR_N  81
`define GTF_COMMON_ADDR_SZ 32
`define GTF_COMMON_DATA_SZ 48

// Attribute addresses
//

`define GTF_COMMON__AEN_QPLL0_FBDIV    32'h00000000
`define GTF_COMMON__AEN_QPLL0_FBDIV_SZ 1

`define GTF_COMMON__AEN_QPLL1_FBDIV    32'h00000001
`define GTF_COMMON__AEN_QPLL1_FBDIV_SZ 1

`define GTF_COMMON__AEN_SDM0TOGGLE    32'h00000002
`define GTF_COMMON__AEN_SDM0TOGGLE_SZ 1

`define GTF_COMMON__AEN_SDM1TOGGLE    32'h00000003
`define GTF_COMMON__AEN_SDM1TOGGLE_SZ 1

`define GTF_COMMON__A_SDM0TOGGLE    32'h00000004
`define GTF_COMMON__A_SDM0TOGGLE_SZ 1

`define GTF_COMMON__A_SDM1DATA_HIGH    32'h00000005
`define GTF_COMMON__A_SDM1DATA_HIGH_SZ 9

`define GTF_COMMON__A_SDM1DATA_LOW    32'h00000006
`define GTF_COMMON__A_SDM1DATA_LOW_SZ 16

`define GTF_COMMON__A_SDM1TOGGLE    32'h00000007
`define GTF_COMMON__A_SDM1TOGGLE_SZ 1

`define GTF_COMMON__BIAS_CFG0    32'h00000008
`define GTF_COMMON__BIAS_CFG0_SZ 16

`define GTF_COMMON__BIAS_CFG1    32'h00000009
`define GTF_COMMON__BIAS_CFG1_SZ 16

`define GTF_COMMON__BIAS_CFG2    32'h0000000a
`define GTF_COMMON__BIAS_CFG2_SZ 16

`define GTF_COMMON__BIAS_CFG3    32'h0000000b
`define GTF_COMMON__BIAS_CFG3_SZ 16

`define GTF_COMMON__BIAS_CFG4    32'h0000000c
`define GTF_COMMON__BIAS_CFG4_SZ 16

`define GTF_COMMON__BIAS_CFG_RSVD    32'h0000000d
`define GTF_COMMON__BIAS_CFG_RSVD_SZ 16

`define GTF_COMMON__COMMON_CFG0    32'h0000000e
`define GTF_COMMON__COMMON_CFG0_SZ 16

`define GTF_COMMON__COMMON_CFG1    32'h0000000f
`define GTF_COMMON__COMMON_CFG1_SZ 16

`define GTF_COMMON__POR_CFG    32'h00000010
`define GTF_COMMON__POR_CFG_SZ 16

`define GTF_COMMON__PPF0_CFG    32'h00000011
`define GTF_COMMON__PPF0_CFG_SZ 16

`define GTF_COMMON__PPF1_CFG    32'h00000012
`define GTF_COMMON__PPF1_CFG_SZ 16

`define GTF_COMMON__QPLL0CLKOUT_RATE    32'h00000013
`define GTF_COMMON__QPLL0CLKOUT_RATE_SZ 32

`define GTF_COMMON__QPLL0_CFG0    32'h00000014
`define GTF_COMMON__QPLL0_CFG0_SZ 16

`define GTF_COMMON__QPLL0_CFG1    32'h00000015
`define GTF_COMMON__QPLL0_CFG1_SZ 16

`define GTF_COMMON__QPLL0_CFG1_G3    32'h00000016
`define GTF_COMMON__QPLL0_CFG1_G3_SZ 16

`define GTF_COMMON__QPLL0_CFG2    32'h00000017
`define GTF_COMMON__QPLL0_CFG2_SZ 16

`define GTF_COMMON__QPLL0_CFG2_G3    32'h00000018
`define GTF_COMMON__QPLL0_CFG2_G3_SZ 16

`define GTF_COMMON__QPLL0_CFG3    32'h00000019
`define GTF_COMMON__QPLL0_CFG3_SZ 16

`define GTF_COMMON__QPLL0_CFG4    32'h0000001a
`define GTF_COMMON__QPLL0_CFG4_SZ 16

`define GTF_COMMON__QPLL0_CP    32'h0000001b
`define GTF_COMMON__QPLL0_CP_SZ 10

`define GTF_COMMON__QPLL0_CP_G3    32'h0000001c
`define GTF_COMMON__QPLL0_CP_G3_SZ 10

`define GTF_COMMON__QPLL0_FBDIV    32'h0000001d
`define GTF_COMMON__QPLL0_FBDIV_SZ 32

`define GTF_COMMON__QPLL0_FBDIV_G3    32'h0000001e
`define GTF_COMMON__QPLL0_FBDIV_G3_SZ 32

`define GTF_COMMON__QPLL0_INIT_CFG0    32'h0000001f
`define GTF_COMMON__QPLL0_INIT_CFG0_SZ 16

`define GTF_COMMON__QPLL0_INIT_CFG1    32'h00000020
`define GTF_COMMON__QPLL0_INIT_CFG1_SZ 8

`define GTF_COMMON__QPLL0_LOCK_CFG    32'h00000021
`define GTF_COMMON__QPLL0_LOCK_CFG_SZ 16

`define GTF_COMMON__QPLL0_LOCK_CFG_G3    32'h00000022
`define GTF_COMMON__QPLL0_LOCK_CFG_G3_SZ 16

`define GTF_COMMON__QPLL0_LPF    32'h00000023
`define GTF_COMMON__QPLL0_LPF_SZ 10

`define GTF_COMMON__QPLL0_LPF_G3    32'h00000024
`define GTF_COMMON__QPLL0_LPF_G3_SZ 10

`define GTF_COMMON__QPLL0_PCI_EN    32'h00000025
`define GTF_COMMON__QPLL0_PCI_EN_SZ 1

`define GTF_COMMON__QPLL0_RATE_SW_USE_DRP    32'h00000026
`define GTF_COMMON__QPLL0_RATE_SW_USE_DRP_SZ 1

`define GTF_COMMON__QPLL0_REFCLK_DIV    32'h00000027
`define GTF_COMMON__QPLL0_REFCLK_DIV_SZ 32

`define GTF_COMMON__QPLL0_SDM_CFG0    32'h00000028
`define GTF_COMMON__QPLL0_SDM_CFG0_SZ 16

`define GTF_COMMON__QPLL0_SDM_CFG1    32'h00000029
`define GTF_COMMON__QPLL0_SDM_CFG1_SZ 16

`define GTF_COMMON__QPLL0_SDM_CFG2    32'h0000002a
`define GTF_COMMON__QPLL0_SDM_CFG2_SZ 16

`define GTF_COMMON__QPLL1CLKOUT_RATE    32'h0000002b
`define GTF_COMMON__QPLL1CLKOUT_RATE_SZ 32

`define GTF_COMMON__QPLL1_CFG0    32'h0000002c
`define GTF_COMMON__QPLL1_CFG0_SZ 16

`define GTF_COMMON__QPLL1_CFG1    32'h0000002d
`define GTF_COMMON__QPLL1_CFG1_SZ 16

`define GTF_COMMON__QPLL1_CFG1_G3    32'h0000002e
`define GTF_COMMON__QPLL1_CFG1_G3_SZ 16

`define GTF_COMMON__QPLL1_CFG2    32'h0000002f
`define GTF_COMMON__QPLL1_CFG2_SZ 16

`define GTF_COMMON__QPLL1_CFG2_G3    32'h00000030
`define GTF_COMMON__QPLL1_CFG2_G3_SZ 16

`define GTF_COMMON__QPLL1_CFG3    32'h00000031
`define GTF_COMMON__QPLL1_CFG3_SZ 16

`define GTF_COMMON__QPLL1_CFG4    32'h00000032
`define GTF_COMMON__QPLL1_CFG4_SZ 16

`define GTF_COMMON__QPLL1_CP    32'h00000033
`define GTF_COMMON__QPLL1_CP_SZ 10

`define GTF_COMMON__QPLL1_CP_G3    32'h00000034
`define GTF_COMMON__QPLL1_CP_G3_SZ 10

`define GTF_COMMON__QPLL1_FBDIV    32'h00000035
`define GTF_COMMON__QPLL1_FBDIV_SZ 32

`define GTF_COMMON__QPLL1_FBDIV_G3    32'h00000036
`define GTF_COMMON__QPLL1_FBDIV_G3_SZ 32

`define GTF_COMMON__QPLL1_INIT_CFG0    32'h00000037
`define GTF_COMMON__QPLL1_INIT_CFG0_SZ 16

`define GTF_COMMON__QPLL1_INIT_CFG1    32'h00000038
`define GTF_COMMON__QPLL1_INIT_CFG1_SZ 8

`define GTF_COMMON__QPLL1_LOCK_CFG    32'h00000039
`define GTF_COMMON__QPLL1_LOCK_CFG_SZ 16

`define GTF_COMMON__QPLL1_LOCK_CFG_G3    32'h0000003a
`define GTF_COMMON__QPLL1_LOCK_CFG_G3_SZ 16

`define GTF_COMMON__QPLL1_LPF    32'h0000003b
`define GTF_COMMON__QPLL1_LPF_SZ 10

`define GTF_COMMON__QPLL1_LPF_G3    32'h0000003c
`define GTF_COMMON__QPLL1_LPF_G3_SZ 10

`define GTF_COMMON__QPLL1_PCI_EN    32'h0000003d
`define GTF_COMMON__QPLL1_PCI_EN_SZ 1

`define GTF_COMMON__QPLL1_RATE_SW_USE_DRP    32'h0000003e
`define GTF_COMMON__QPLL1_RATE_SW_USE_DRP_SZ 1

`define GTF_COMMON__QPLL1_REFCLK_DIV    32'h0000003f
`define GTF_COMMON__QPLL1_REFCLK_DIV_SZ 32

`define GTF_COMMON__QPLL1_SDM_CFG0    32'h00000040
`define GTF_COMMON__QPLL1_SDM_CFG0_SZ 16

`define GTF_COMMON__QPLL1_SDM_CFG1    32'h00000041
`define GTF_COMMON__QPLL1_SDM_CFG1_SZ 16

`define GTF_COMMON__QPLL1_SDM_CFG2    32'h00000042
`define GTF_COMMON__QPLL1_SDM_CFG2_SZ 16

`define GTF_COMMON__RSVD_ATTR0    32'h00000043
`define GTF_COMMON__RSVD_ATTR0_SZ 16

`define GTF_COMMON__RSVD_ATTR1    32'h00000044
`define GTF_COMMON__RSVD_ATTR1_SZ 16

`define GTF_COMMON__RSVD_ATTR2    32'h00000045
`define GTF_COMMON__RSVD_ATTR2_SZ 16

`define GTF_COMMON__RSVD_ATTR3    32'h00000046
`define GTF_COMMON__RSVD_ATTR3_SZ 16

`define GTF_COMMON__RXRECCLKOUT0_SEL    32'h00000047
`define GTF_COMMON__RXRECCLKOUT0_SEL_SZ 2

`define GTF_COMMON__RXRECCLKOUT1_SEL    32'h00000048
`define GTF_COMMON__RXRECCLKOUT1_SEL_SZ 2

`define GTF_COMMON__SARC_ENB    32'h00000049
`define GTF_COMMON__SARC_ENB_SZ 1

`define GTF_COMMON__SARC_SEL    32'h0000004a
`define GTF_COMMON__SARC_SEL_SZ 1

`define GTF_COMMON__SDM0INITSEED0_0    32'h0000004b
`define GTF_COMMON__SDM0INITSEED0_0_SZ 16

`define GTF_COMMON__SDM0INITSEED0_1    32'h0000004c
`define GTF_COMMON__SDM0INITSEED0_1_SZ 9

`define GTF_COMMON__SDM1INITSEED0_0    32'h0000004d
`define GTF_COMMON__SDM1INITSEED0_0_SZ 16

`define GTF_COMMON__SDM1INITSEED0_1    32'h0000004e
`define GTF_COMMON__SDM1INITSEED0_1_SZ 9

`define GTF_COMMON__SIM_MODE    32'h0000004f
`define GTF_COMMON__SIM_MODE_SZ 48

`define GTF_COMMON__SIM_RESET_SPEEDUP    32'h00000050
`define GTF_COMMON__SIM_RESET_SPEEDUP_SZ 40

`endif  // B_GTF_COMMON_DEFINES_VH