`include "B_IBUFDS_IBUFDISABLE_INT_defines.vh"

reg [`IBUFDS_IBUFDISABLE_INT_DATA_SZ-1:0] ATTR [0:`IBUFDS_IBUFDISABLE_INT_ADDR_N-1];
reg [`IBUFDS_IBUFDISABLE_INT__DIFF_TERM_SZ:1] DIFF_TERM_REG = DIFF_TERM;
reg [`IBUFDS_IBUFDISABLE_INT__DQS_BIAS_SZ:1] DQS_BIAS_REG = DQS_BIAS;
reg [`IBUFDS_IBUFDISABLE_INT__IBUF_LOW_PWR_SZ:1] IBUF_LOW_PWR_REG = IBUF_LOW_PWR;
reg [`IBUFDS_IBUFDISABLE_INT__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IBUFDS_IBUFDISABLE_INT__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IBUFDS_IBUFDISABLE_INT__DIFF_TERM] = DIFF_TERM;
  ATTR[`IBUFDS_IBUFDISABLE_INT__DQS_BIAS] = DQS_BIAS;
  ATTR[`IBUFDS_IBUFDISABLE_INT__IBUF_LOW_PWR] = IBUF_LOW_PWR;
  ATTR[`IBUFDS_IBUFDISABLE_INT__IOSTANDARD] = IOSTANDARD;
  ATTR[`IBUFDS_IBUFDISABLE_INT__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  DIFF_TERM_REG = ATTR[`IBUFDS_IBUFDISABLE_INT__DIFF_TERM];
  DQS_BIAS_REG = ATTR[`IBUFDS_IBUFDISABLE_INT__DQS_BIAS];
  IBUF_LOW_PWR_REG = ATTR[`IBUFDS_IBUFDISABLE_INT__IBUF_LOW_PWR];
  IOSTANDARD_REG = ATTR[`IBUFDS_IBUFDISABLE_INT__IOSTANDARD];
  USE_IBUFDISABLE_REG = ATTR[`IBUFDS_IBUFDISABLE_INT__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IBUFDS_IBUFDISABLE_INT_ADDR_SZ-1:0] addr;
  input  [`IBUFDS_IBUFDISABLE_INT_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IBUFDS_IBUFDISABLE_INT_DATA_SZ-1:0] read_attr;
  input  [`IBUFDS_IBUFDISABLE_INT_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
