----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description : This module implement the parallel loopback function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
use phy_plus_lane_lib.all;

entity parallel_loopback is
   port (
      CLK                              : in  std_logic;                          --! Clock generated by GTY IP
      RST_N                            : in  std_logic;                          --! Global reset
      -- FROM lane_ctrl_word_insert
      DATA_TX_FROM_LCWI                : in  std_logic_vector(31 downto 00);     --! 32-bit Data
      VALID_K_CARAC_FROM_LCWI          : in  std_logic_vector(03 downto 00);     --! 4-bit Valid K character
      DATA_RDY_FROM_LCWI               : in  std_logic;                          --! Data ready flag
      -- FROM rx_sync_fsm
      DATA_TX_FROM_RSF                 : in  std_logic_vector(31 downto 00);     --! 32-bit Data
      VALID_K_CARAC_FROM_RSF           : in  std_logic_vector(03 downto 00);     --! 4-bit Valid K character
      DATA_RDY_FROM_RSF                : in  std_logic;                          --! Data ready flag
      --FROM skip_insertion
      WAIT_SKIP_DATA                   : in  std_logic;                          --! Wait for data to be skip
      --TO lane_ctrl_word_detection
      DATA_TX_TO_LCWD                  : out std_logic_vector(31 downto 00);     --! 32-bit Data
      VALID_K_CARAC_TO_LCWD            : out std_logic_vector(03 downto 00);     --! 4-bit Valid K character
      DATA_RDY_TO_LCWD                 : out std_logic;                          --! Data ready flag
      -- Parameter
      PARALLEL_LOOPBACK_EN             : in  std_logic                           --! Enable or disable the parallel loopback for the lane
   );
end parallel_loopback;

architecture rtl of parallel_loopback is
----------------------------- Declaration signals -----------------------------
signal wait_skip_data_r                : std_logic;                              --! 
signal wait_skip_data_rr               : std_logic;
signal wait_skip_data_rrr              : std_logic;

begin
   p_delay_wait_skip : process(CLK, RST_N)
   begin
      if RST_N = '0' then
         wait_skip_data_r   <= '0';
         wait_skip_data_rr  <= '0';
         wait_skip_data_rrr <= '0';
      elsif rising_edge(CLK) then
         wait_skip_data_r      <= WAIT_SKIP_DATA;
         wait_skip_data_rr     <= wait_skip_data_r;
         wait_skip_data_rrr    <= wait_skip_data_rr;
      end if;
   end process p_delay_wait_skip;
   
   -- Allows to make a parallele loopback into the LANE layer
   DATA_TX_TO_LCWD       <= DATA_TX_FROM_LCWI       when PARALLEL_LOOPBACK_EN = '1' else DATA_TX_FROM_RSF;
   VALID_K_CARAC_TO_LCWD <= VALID_K_CARAC_FROM_LCWI when PARALLEL_LOOPBACK_EN = '1' else VALID_K_CARAC_FROM_RSF;
   DATA_RDY_TO_LCWD      <= (DATA_RDY_FROM_LCWI and not(wait_skip_data_rrr) )    when PARALLEL_LOOPBACK_EN = '1' else DATA_RDY_FROM_RSF;

end architecture rtl;