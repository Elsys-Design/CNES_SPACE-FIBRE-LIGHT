`include "B_DSP_FPM_PIPEREG_TEST_defines.vh"

reg [`DSP_FPM_PIPEREG_TEST_DATA_SZ-1:0] ATTR [0:`DSP_FPM_PIPEREG_TEST_ADDR_N-1];
reg [24:1] A_FPTYPE_REG = A_FPTYPE;
reg [24:1] B_D_FPTYPE_REG = B_D_FPTYPE;
reg [56:1] EN_SCAN_REG = EN_SCAN;
reg [31:0] FPMPIPEREG_REG = FPMPIPEREG;
reg IS_RSTFPMPIPE_INVERTED_REG = IS_RSTFPMPIPE_INVERTED;
reg [40:1] LEGACY_REG = LEGACY;
reg [31:0] MREG_REG = MREG;
reg [40:1] RESET_MODE_REG = RESET_MODE;
reg [64:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_FPM_PIPEREG_TEST__A_FPTYPE] = A_FPTYPE;
  ATTR[`DSP_FPM_PIPEREG_TEST__B_D_FPTYPE] = B_D_FPTYPE;
  ATTR[`DSP_FPM_PIPEREG_TEST__EN_SCAN] = EN_SCAN;
  ATTR[`DSP_FPM_PIPEREG_TEST__FPMPIPEREG] = FPMPIPEREG;
  ATTR[`DSP_FPM_PIPEREG_TEST__IS_RSTFPMPIPE_INVERTED] = IS_RSTFPMPIPE_INVERTED;
  ATTR[`DSP_FPM_PIPEREG_TEST__LEGACY] = LEGACY;
  ATTR[`DSP_FPM_PIPEREG_TEST__MREG] = MREG;
  ATTR[`DSP_FPM_PIPEREG_TEST__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_FPM_PIPEREG_TEST__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  A_FPTYPE_REG = ATTR[`DSP_FPM_PIPEREG_TEST__A_FPTYPE];
  B_D_FPTYPE_REG = ATTR[`DSP_FPM_PIPEREG_TEST__B_D_FPTYPE];
  EN_SCAN_REG = ATTR[`DSP_FPM_PIPEREG_TEST__EN_SCAN];
  FPMPIPEREG_REG = ATTR[`DSP_FPM_PIPEREG_TEST__FPMPIPEREG];
  IS_RSTFPMPIPE_INVERTED_REG = ATTR[`DSP_FPM_PIPEREG_TEST__IS_RSTFPMPIPE_INVERTED];
  LEGACY_REG = ATTR[`DSP_FPM_PIPEREG_TEST__LEGACY];
  MREG_REG = ATTR[`DSP_FPM_PIPEREG_TEST__MREG];
  RESET_MODE_REG = ATTR[`DSP_FPM_PIPEREG_TEST__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_FPM_PIPEREG_TEST__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FPM_PIPEREG_TEST_ADDR_SZ-1:0] addr;
  input  [`DSP_FPM_PIPEREG_TEST_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FPM_PIPEREG_TEST_DATA_SZ-1:0] read_attr;
  input  [`DSP_FPM_PIPEREG_TEST_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
