----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module describe the Output Buffer & Flow control
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_link_reset is
  port (
    RST_N                   : in  std_logic;                                    --! global reset
    CLK                     : in  std_logic;                                    --! Clock generated by GTY IP
    -- Link Reset
    LINK_RESET_DLRE         : out std_logic;
    -- Lane interface
    LANE_RESET_DLRE         : out std_logic;
    --MIB interface
    INTERFACE_RESET_MIB     : in std_logic;
    LINK_RESET_MIB              : in std_logic;

  );
end data_link_reset;

architecture rtl of data_link_reset is
----------------------------- Declaration signals -----------------------------
  type link_rst_fsm is (
    CONF_RST_ST,
    NEAR_END_RST_ST,
    CHECK_FAR_END_RST_ST,
    LINK_INIT_ST
  );

  signal current_state          : link_rst_fsm;
  signal current_state_fct      : req_fct_fsm; 

begin
---------------------------------------------------------
-----                     Assignation               -----
---------------------------------------------------------
---------------------------------------------------------
-----                     Instanciation             -----
---------------------------------------------------------
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------

---------------------------------------------------------
-- Process: p_data_in_fifo
-- Description: Manages the data written into the fifo
---------------------------------------------------------
p_data_in_fifo: process(CLK, RST_N)
begin
  if RST_N = '0' then
    current_state   <= CONF_RST_ST;
    LINK_RESET_DLRE <= '0';
    LANE_RESET_DLRE <= '0';
  elsif rising_edge(CLK) then
    case current_state is 
      when CONF_RST_ST          =>
                                  LINK_RESET_DLRE <= '1';
                                  LANE_RESET_DLRE <= '1';
                                  current_state   <= CONF_RST_ST;
      when NEAR_END_RST_ST      => 
                                  LINK_RESET_DLRE <= '1';
                                  LANE_RESET_DLRE <= '1';
                                  if INTERFACE_RESET_MIB ='1' then
                                    current_state   <= CONF_RST_ST;
                                  else
                                    current_state   <= CHECK_FAR_END_RST_ST;
                                  end if;
      when CHECK_FAR_END_RST_ST => 
                                  if INTERFACE_RESET_MIB ='1' then
                                    current_state   <= CONF_RST_ST;
                                  elsif LINK_RESET_MIB  ='1' then 
                                    current_state   <= NEAR_END_RST_ST;
                                  end if;
      when LINK_INIT_ST         => 
                                  if INTERFACE_RESET_MIB ='1' then
                                    current_state   <= CONF_RST_ST;
                                  elsif LINK_RESET_MIB  ='1' then 
                                    current_state   <= NEAR_END_RST_ST;
                                  end if;
    end case;
  end if;
end process p_data_in_fifo;
end architecture rtl;