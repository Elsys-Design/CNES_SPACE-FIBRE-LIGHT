// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_PREADD_DATA_DEFINES_VH
`else
`define B_DSP_PREADD_DATA_DEFINES_VH

// Look-up table parameters
//

`define DSP_PREADD_DATA_ADDR_N  11
`define DSP_PREADD_DATA_ADDR_SZ 32
`define DSP_PREADD_DATA_DATA_SZ 64

// Attribute addresses
//

`define DSP_PREADD_DATA__ADREG    32'h00000000
`define DSP_PREADD_DATA__ADREG_SZ 32

`define DSP_PREADD_DATA__AMULTSEL    32'h00000001
`define DSP_PREADD_DATA__AMULTSEL_SZ 16

`define DSP_PREADD_DATA__BMULTSEL    32'h00000002
`define DSP_PREADD_DATA__BMULTSEL_SZ 16

`define DSP_PREADD_DATA__DREG    32'h00000003
`define DSP_PREADD_DATA__DREG_SZ 32

`define DSP_PREADD_DATA__INMODEREG    32'h00000004
`define DSP_PREADD_DATA__INMODEREG_SZ 32

`define DSP_PREADD_DATA__IS_CLK_INVERTED    32'h00000005
`define DSP_PREADD_DATA__IS_CLK_INVERTED_SZ 1

`define DSP_PREADD_DATA__IS_INMODE_INVERTED    32'h00000006
`define DSP_PREADD_DATA__IS_INMODE_INVERTED_SZ 5

`define DSP_PREADD_DATA__IS_RSTD_INVERTED    32'h00000007
`define DSP_PREADD_DATA__IS_RSTD_INVERTED_SZ 1

`define DSP_PREADD_DATA__IS_RSTINMODE_INVERTED    32'h00000008
`define DSP_PREADD_DATA__IS_RSTINMODE_INVERTED_SZ 1

`define DSP_PREADD_DATA__PREADDINSEL    32'h00000009
`define DSP_PREADD_DATA__PREADDINSEL_SZ 8

`define DSP_PREADD_DATA__USE_MULT    32'h0000000a
`define DSP_PREADD_DATA__USE_MULT_SZ 64

`endif  // B_DSP_PREADD_DATA_DEFINES_VH