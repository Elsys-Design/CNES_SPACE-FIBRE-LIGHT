// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_PREADD_DATA58_DEFINES_VH
`else
`define B_DSP_PREADD_DATA58_DEFINES_VH

// Look-up table parameters
//

`define DSP_PREADD_DATA58_ADDR_N  16
`define DSP_PREADD_DATA58_ADDR_SZ 32
`define DSP_PREADD_DATA58_DATA_SZ 64

// Attribute addresses
//

`define DSP_PREADD_DATA58__ADREG    32'h00000000
`define DSP_PREADD_DATA58__ADREG_SZ 32

`define DSP_PREADD_DATA58__AMULTSEL    32'h00000001
`define DSP_PREADD_DATA58__AMULTSEL_SZ 16

`define DSP_PREADD_DATA58__AREG    32'h00000002
`define DSP_PREADD_DATA58__AREG_SZ 32

`define DSP_PREADD_DATA58__BMULTSEL    32'h00000003
`define DSP_PREADD_DATA58__BMULTSEL_SZ 16

`define DSP_PREADD_DATA58__BREG    32'h00000004
`define DSP_PREADD_DATA58__BREG_SZ 32

`define DSP_PREADD_DATA58__DREG    32'h00000005
`define DSP_PREADD_DATA58__DREG_SZ 32

`define DSP_PREADD_DATA58__DSP_MODE    32'h00000006
`define DSP_PREADD_DATA58__DSP_MODE_SZ 48

`define DSP_PREADD_DATA58__INMODEREG    32'h00000007
`define DSP_PREADD_DATA58__INMODEREG_SZ 32

`define DSP_PREADD_DATA58__IS_INMODE_INVERTED    32'h00000008
`define DSP_PREADD_DATA58__IS_INMODE_INVERTED_SZ 5

`define DSP_PREADD_DATA58__IS_NEGATE_INVERTED    32'h00000009
`define DSP_PREADD_DATA58__IS_NEGATE_INVERTED_SZ 3

`define DSP_PREADD_DATA58__IS_RSTINMODE_INVERTED    32'h0000000a
`define DSP_PREADD_DATA58__IS_RSTINMODE_INVERTED_SZ 1

`define DSP_PREADD_DATA58__LEGACY    32'h0000000b
`define DSP_PREADD_DATA58__LEGACY_SZ 40

`define DSP_PREADD_DATA58__MREG    32'h0000000c
`define DSP_PREADD_DATA58__MREG_SZ 32

`define DSP_PREADD_DATA58__PREADDINSEL    32'h0000000d
`define DSP_PREADD_DATA58__PREADDINSEL_SZ 8

`define DSP_PREADD_DATA58__RESET_MODE    32'h0000000e
`define DSP_PREADD_DATA58__RESET_MODE_SZ 40

`define DSP_PREADD_DATA58__USE_MULT    32'h0000000f
`define DSP_PREADD_DATA58__USE_MULT_SZ 64

`endif  // B_DSP_PREADD_DATA58_DEFINES_VH