-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 17/07/2025
--
-- Description : This is the testbench of the ppl_64_lane_ctrl_word_insert module  
----------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library work;
   use work.pkg_simu.all;

entity tb_ppl_64_lane_ctrl_word_insert is
end entity;

architecture tb of tb_ppl_64_lane_ctrl_word_insert is

component ppl_64_lane_ctrl_word_insert is
  port (
    RST_N                                : in  std_logic;                                          --! global reset
    CLK                                  : in  std_logic;                                          --! Clock generated by HSSL IP
    -- Data-Link interface
    RD_DATA_EN_PLCWI                           : out std_logic;                                          --! Read command to receive data from Data-link layer
    RD_DATA_VALID_DL                     : in  std_logic;                                          --! Data valid flag from Data-link layer
    CAPABILITY_DL                        : in  std_logic_vector(7 downto 0);                       --! Capability field from DATA-LINK layer
    DATA_TX_DL                           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit receive from DATA_LINK layer
    VALID_K_CHARAC_DL                    : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character from DATA-LINK layer
    NO_DATA_DL                           : in  std_logic;                                          --! Flag to enable the send of IDLE words when no data should be available from Data-Link
    -- ppl_64_skip_insertion (PLSI) interface
    WAIT_SEND_DATA_PLSI                  : in  std_logic;                                          --! Flag to indicates that the skip_insertion send a SKIP control word
    NEW_DATA_PLCWI                       : out std_logic;                                          --! New data send to skip_insertion
    DATA_TX_PLCWI                        : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit send to manufacturer IP
    VALID_K_CHARAC_PLCWI                 : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character
    -- ppl_64_lane_init_fsm (PLIF) interface
    SEND_INIT1_CTRL_WORD_PLIF           : in  std_logic;                                          --! Flag to send INIT1 control word following by 64 pseudo-random data words
    SEND_INIT2_CTRL_WORD_PLIF           : in  std_logic;                                          --! Flag to send INIT2 control word following by 64 pseudo-random data words
    SEND_INIT3_CTRL_WORD_PLIF           : in  std_logic;                                          --! Flag to send INIT3 control word following by 64 pseudo-random data words
    ENABLE_TRANSM_DATA_PLIF             : in  std_logic;                                          --! Flag to enable to send data
    SEND_32_STANDBY_CTRL_WORDS_PLIF     : in  std_logic;                                          --! Flag to send STANDBY control word x32
    SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF : in  std_logic;                                          --! Flag to send LOSS_SIGNAL control word x32
    STANDBY_SIGNAL_X32_PLCWI             : out std_logic;                                          --! Flag STANDBY control word has been send x32
    LOST_SIGNAL_X32_PLCWI                : out std_logic;                                          --! Flag LOST_SIGNAL control word has been send x32
    -- MIB interface
    STANDBY_REASON_MIB                   : in  std_logic_vector(7 downto 0);                       --! Standby reason from MIB
    LOST_CAUSE_MIB                       : in  std_logic_vector(1 downto 0)                        --! Flag to indicate the reason of the LOST_SIGNAL
  );
end component;


---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
constant periode                              : time := 13.334 ns;

signal RST_N                                  : std_logic := '0';
signal CLK                                    : std_logic := '0';

signal RD_DATA_EN_PLCWI                             : std_logic;
signal RD_DATA_VALID_DL                       : std_logic:='0';
signal CAPABILITY_DL                          : std_logic_vector(7 downto 0) := (others => '0');
signal DATA_TX_DL                             : std_logic_vector(C_DATA_LENGTH-1 downto 0) := (others => '0');
signal VALID_K_CHARAC_DL                      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0) := (others => '0');
signal NO_DATA_DL                             : std_logic := '0';
signal WAIT_SEND_DATA_PLSI                    : std_logic := '0';
signal NEW_DATA_PLCWI                         : std_logic;
signal DATA_TX_PLCWI                          : std_logic_vector(C_DATA_LENGTH-1 downto 0);
signal VALID_K_CHARAC_PLCWI                   : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
signal SEND_INIT1_CTRL_WORD_PLIF             : std_logic := '0';
signal SEND_INIT2_CTRL_WORD_PLIF             : std_logic := '0';
signal SEND_INIT3_CTRL_WORD_PLIF             : std_logic := '0';
signal ENABLE_TRANSM_DATA_PLIF               : std_logic := '0';
signal SEND_32_STANDBY_CTRL_WORDS_PLIF       : std_logic := '0';
signal STANDBY_REASON_MIB                     : std_logic_vector(7 downto 0) := (others => '0');
signal SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF   : std_logic := '0';
signal LOST_CAUSE_MIB                         : std_logic_vector(1 downto 0) := (others => '0');
signal STANDBY_SIGNAL_X32_PLCWI               : std_logic;
signal LOST_SIGNAL_X32_PLCWI                  : std_logic;

begin

---------------------------------------------------------
-----                  Instantiation                -----
---------------------------------------------------------
DUT : ppl_64_lane_ctrl_word_insert
port map(
   RST_N                                => RST_N,
   CLK                                  => CLK,
   RD_DATA_EN_PLCWI                           => RD_DATA_EN_PLCWI,
   RD_DATA_VALID_DL                     => RD_DATA_VALID_DL,
   CAPABILITY_DL                        => CAPABILITY_DL,
   DATA_TX_DL                           => DATA_TX_DL,
   VALID_K_CHARAC_DL                    => VALID_K_CHARAC_DL,
   NO_DATA_DL                           => NO_DATA_DL,
   WAIT_SEND_DATA_PLSI                  => WAIT_SEND_DATA_PLSI ,
   NEW_DATA_PLCWI                       => NEW_DATA_PLCWI,
   DATA_TX_PLCWI                        => DATA_TX_PLCWI,
   VALID_K_CHARAC_PLCWI                 => VALID_K_CHARAC_PLCWI,
   SEND_INIT1_CTRL_WORD_PLIF           => SEND_INIT1_CTRL_WORD_PLIF,
   SEND_INIT2_CTRL_WORD_PLIF           => SEND_INIT2_CTRL_WORD_PLIF,
   SEND_INIT3_CTRL_WORD_PLIF           => SEND_INIT3_CTRL_WORD_PLIF,
   ENABLE_TRANSM_DATA_PLIF             => ENABLE_TRANSM_DATA_PLIF,
   SEND_32_STANDBY_CTRL_WORDS_PLIF     => SEND_32_STANDBY_CTRL_WORDS_PLIF,
   SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF => SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF,
   STANDBY_SIGNAL_X32_PLCWI             => STANDBY_SIGNAL_X32_PLCWI,
   LOST_SIGNAL_X32_PLCWI                => LOST_SIGNAL_X32_PLCWI,
   STANDBY_REASON_MIB                   => STANDBY_REASON_MIB,
   LOST_CAUSE_MIB                       => LOST_CAUSE_MIB
);

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
-- generate clock 150 MHz
horloge : process
begin
   CLK   <= not CLK;
   wait for periode/2;
end process;

scenario : process
   variable test_failed : boolean := false;
begin
  RST_N <= '0';
  wait for 10 us;
  wait until rising_edge(CLK);
  RST_N <= '1';
  wait for 20 us;

  --------------------------------------
  -- TEST 0: INIT Control Word        --
  --------------------------------------
  -- Test 0: INIT 1
  --------------------------------------
  SEND_INIT1_CTRL_WORD_PLIF <= '1';
  wait until rising_edge(CLK) and NEW_DATA_PLCWI ='1';
  for i in 0 to 31 loop
    check_equal("Test 0: INIT 1: DATA_TX_PLCWI i="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2+1,32))& std_logic_vector(to_unsigned(i*2,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 1: VALID_K_CHARAC_PLCWI i="& integer'image(i), x"00",                                                                          VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 1: NEW_DATA_PLCWI i="& integer'image(i),       '1',                                                                            NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 1 on word 0
  check_equal("Test 0: INIT 1: DATA_TX_PLCWI i=C_INIT1_WORD word 0"     ,    std_logic_vector(to_unsigned(0,32)) & C_INIT1_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 1: VALID_K_CHARAC_PLCWI i= C_INIT1_WORD word 0", x"01",                                              VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 1: NEW_DATA_PLCWI i= C_INIT1_WORD word 0",       '1',                                                NEW_DATA_PLCWI,       test_failed);
  wait until rising_edge(CLK);
  for i in 1 to 31 loop
    check_equal("Test 0: INIT 1: DATA_TX_PLCWI i2="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2,32))& std_logic_vector(to_unsigned((i-1)*2+1,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 1: VALID_K_CHARAC_PLCWI i2="& integer'image(i), x"00",                                                                              VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 1: NEW_DATA_PLCWI i2="& integer'image(i),       '1',                                                                                NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 1 on word 1
  check_equal("Test 0: INIT 1: DATA_TX_PLCWI i=C_INIT1_WORD word 1"     ,    C_INIT1_WORD & std_logic_vector(to_unsigned(63,32)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 1: VALID_K_CHARAC_PLCWI i= C_INIT1_WORD word 1", x"10",                                               VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 1: NEW_DATA_PLCWI i= C_INIT1_WORD word 1",       '1',                                                 NEW_DATA_PLCWI,       test_failed);
  SEND_INIT1_CTRL_WORD_PLIF <= '0';
  wait for 10 us;
  -- Test 0: INIT 2
  --------------------------------------
  wait until falling_edge(CLK);
  SEND_INIT2_CTRL_WORD_PLIF <= '1';
  wait until rising_edge(CLK) and NEW_DATA_PLCWI ='1';
  for i in 0 to 31 loop
    check_equal("Test 0: INIT 2: DATA_TX_PLCWI i="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2+1,32))& std_logic_vector(to_unsigned(i*2,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 2: VALID_K_CHARAC_PLCWI i="& integer'image(i), x"00",                                                                          VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 2: NEW_DATA_PLCWI i="& integer'image(i),       '1',                                                                            NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 2 on word 0
  check_equal("Test 0: INIT 2: DATA_TX_PLCWI i=C_INIT2_WORD word 0"     ,    std_logic_vector(to_unsigned(0,32)) & C_INIT2_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 2: VALID_K_CHARAC_PLCWI i= C_INIT2_WORD word 0", x"01",                                              VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 2: NEW_DATA_PLCWI i= C_INIT2_WORD word 0",       '1',                                                NEW_DATA_PLCWI,       test_failed);
  wait until rising_edge(CLK);
  for i in 1 to 31 loop
    check_equal("Test 0: INIT 2: DATA_TX_PLCWI i2="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2,32))& std_logic_vector(to_unsigned((i-1)*2+1,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 2: VALID_K_CHARAC_PLCWI i2="& integer'image(i), x"00",                                                                              VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 2: NEW_DATA_PLCWI i2="& integer'image(i),       '1',                                                                                NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 2 on word 1
  check_equal("Test 0: INIT 2: DATA_TX_PLCWI i=C_INIT2_WORD word 1"     ,    C_INIT2_WORD & std_logic_vector(to_unsigned(63,32)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 2: VALID_K_CHARAC_PLCWI i= C_INIT2_WORD word 1", x"10",                                               VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 2: NEW_DATA_PLCWI i= C_INIT2_WORD word 1",       '1',                                                 NEW_DATA_PLCWI,       test_failed);
  SEND_INIT2_CTRL_WORD_PLIF <= '0';
  wait for 10 us;
  -- Test 0: INIT 3
  --------------------------------------
  wait until falling_edge(CLK);
  SEND_INIT3_CTRL_WORD_PLIF <= '1';
  CAPABILITY_DL  <= x"FF";
  wait until rising_edge(CLK) and NEW_DATA_PLCWI ='1';
  for i in 0 to 31 loop
    check_equal("Test 0: INIT 3: DATA_TX_PLCWI i="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2+1,32))& std_logic_vector(to_unsigned(i*2,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 3: VALID_K_CHARAC_PLCWI i="& integer'image(i), x"00",                                                                          VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 3: NEW_DATA_PLCWI i="& integer'image(i),       '1',                                                                            NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 3 on word 0
  check_equal("Test 0: INIT 3: DATA_TX_PLCWI i=C_INIT3_WORD word 0"     ,    std_logic_vector(to_unsigned(0,32)) & x"FF" & C_INIT3_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 3: VALID_K_CHARAC_PLCWI i= C_INIT3_WORD word 0", x"01",                                                      VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 3: NEW_DATA_PLCWI i= C_INIT3_WORD word 0",       '1',                                                        NEW_DATA_PLCWI,       test_failed);
  wait until rising_edge(CLK);
  for i in 1 to 31 loop
    check_equal("Test 0: INIT 3: DATA_TX_PLCWI i2="& integer'image(i)    ,    std_logic_vector(to_unsigned(i*2,32))& std_logic_vector(to_unsigned((i-1)*2+1,32)), DATA_TX_PLCWI,        test_failed);
    check_equal("Test 0: INIT 3: VALID_K_CHARAC_PLCWI i2="& integer'image(i), x"00",                                                                              VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 0: INIT 3: NEW_DATA_PLCWI i2="& integer'image(i),       '1',                                                                                NEW_DATA_PLCWI,       test_failed);
    wait until rising_edge(CLK);
  end loop;
  -- Check INIT 3 on word 1
  check_equal("Test 0: INIT 3: DATA_TX_PLCWI i=C_INIT3_WORD word 1"     ,    x"FF" & C_INIT3_WORD & std_logic_vector(to_unsigned(63,32)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 0: INIT 3: VALID_K_CHARAC_PLCWI i= C_INIT3_WORD word 1", x"10",                                                       VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 0: INIT 3: NEW_DATA_PLCWI i= C_INIT3_WORD word 1",       '1',                                                         NEW_DATA_PLCWI,       test_failed);
  SEND_INIT3_CTRL_WORD_PLIF <= '0';
  -----------------------------------------
  -- TEST 1: Active state: transmit Data --
  -----------------------------------------
  NO_DATA_DL           <= '1';
  wait for 10 us;
  wait until falling_edge(CLK);
  -- Tests active_st no data from DL
  ENABLE_TRANSM_DATA_PLIF   <= '1';
  wait until falling_edge(CLK);
  check_equal("Test 1: No data dl: DATA_TX_PLCWI"     ,   C_IDLE_WORD & C_IDLE_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: No data dl: VALID_K_CHARAC_PLCWI", x"11",                     VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: No data dl: NEW_DATA_PLCWI",       '1' ,                      NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: No data dl: RD_DATA_EN_PLCWI",           '1' ,                      RD_DATA_EN_PLCWI,           test_failed);
  -- Test active state with data
  NO_DATA_DL           <= '0';
  RD_DATA_VALID_DL     <= '1';
  DATA_TX_DL           <= std_logic_vector(to_unsigned(1,DATA_TX_DL'length));
  VALID_K_CHARAC_DL    <= x"00";
  wait until falling_edge(CLK);
  check_equal("Test 1: transmit data: DATA_TX_PLCWI"     ,   std_logic_vector(to_unsigned(1,DATA_TX_DL'length)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: transmit data: VALID_K_CHARAC_PLCWI", x"00",                                              VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: transmit data: NEW_DATA_PLCWI",       '1' ,                                               NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: transmit data: RD_DATA_EN_PLCWI",           '1' ,                                               RD_DATA_EN_PLCWI,           test_failed);

  DATA_TX_DL           <= std_logic_vector(to_unsigned(200,DATA_TX_DL'length));
  VALID_K_CHARAC_DL    <= x"00";
  wait until falling_edge(CLK);
  check_equal("Test 1: transmit data: DATA_TX_PLCWI"     ,   std_logic_vector(to_unsigned(200,DATA_TX_DL'length)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: transmit data: VALID_K_CHARAC_PLCWI", x"00",                                                VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: transmit data: NEW_DATA_PLCWI",       '1' ,                                                 NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: transmit data: RD_DATA_EN_PLCWI",           '1' ,                                                 RD_DATA_EN_PLCWI,           test_failed);
  -- No RD DATA VALID
  RD_DATA_VALID_DL     <= '0';
  wait until falling_edge(CLK);
  check_equal("Test 1: No RD DATA VALID: DATA_TX_PLCWI"     ,   C_IDLE_WORD & C_IDLE_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: No RD DATA VALID: VALID_K_CHARAC_PLCWI", x"11",                     VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: No RD DATA VALID: NEW_DATA_PLCWI",       '1' ,                      NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: No RD DATA VALID: RD_DATA_EN_PLCWI",           '1' ,                      RD_DATA_EN_PLCWI,           test_failed);
  -- WAIT_SEND_DATA_PLSI at '1'
  WAIT_SEND_DATA_PLSI  <= '1';
  RD_DATA_VALID_DL     <= '1';
  wait until falling_edge(CLK);
  check_equal("Test 1: WAIT_SEND_DATA_PLSI: DATA_TX_PLCWI"     ,   std_logic_vector(to_unsigned(200,DATA_TX_DL'length)), DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: WAIT_SEND_DATA_PLSI: VALID_K_CHARAC_PLCWI", x"00",                                                VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: WAIT_SEND_DATA_PLSI: NEW_DATA_PLCWI",       '1' ,                                                 NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: WAIT_SEND_DATA_PLSI: RD_DATA_EN_PLCWI",           '0' ,                                                 RD_DATA_EN_PLCWI,           test_failed);

  RD_DATA_VALID_DL     <= '0';
  wait until falling_edge(CLK);
  check_equal("Test 1: WAIT_SEND_DATA_PLSI: DATA_TX_PLCWI"     ,   C_IDLE_WORD & C_IDLE_WORD, DATA_TX_PLCWI,        test_failed);
  check_equal("Test 1: WAIT_SEND_DATA_PLSI: VALID_K_CHARAC_PLCWI", x"11",                     VALID_K_CHARAC_PLCWI, test_failed);
  check      ("Test 1: WAIT_SEND_DATA_PLSI: NEW_DATA_PLCWI",       '1' ,                      NEW_DATA_PLCWI,       test_failed);
  check      ("Test 1: WAIT_SEND_DATA_PLSI: RD_DATA_EN_PLCWI",           '0' ,                      RD_DATA_EN_PLCWI,           test_failed);
  ENABLE_TRANSM_DATA_PLIF   <= '0';
  wait for 10 us;
  --------------------------------------
  -- TEST 2:  Standby Control Word    --
  --------------------------------------
  -- test STANDBY
  SEND_32_STANDBY_CTRL_WORDS_PLIF <= '1';
  STANDBY_REASON_MIB             <= x"FF";
  wait until falling_edge(CLK);
  for i in 0 to 15 loop
    wait until falling_edge(CLK);
    check_equal("Test 2: Standby Control Word: DATA_TX_PLCWI i="& integer'image(i)    ,    x"FF" & C_STANDBY_WORD & x"FF" & C_STANDBY_WORD, DATA_TX_PLCWI,        test_failed);
    check_equal("Test 2: Standby Control Word: VALID_K_CHARAC_PLCWI i="& integer'image(i), x"11",                                           VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 2: Standby Control Word: NEW_DATA_PLCWI i="& integer'image(i),       '1' ,                                            NEW_DATA_PLCWI,       test_failed);
    check      ("Test 2: Standby Control Word: STANDBY_SIGNAL_X32_PLCWI i="& integer'image(i),   '0' ,                                            STANDBY_SIGNAL_X32_PLCWI,   test_failed);
  end loop;
  wait until falling_edge(CLK);
  check      ("Test 2: Standby Control Word: STANDBY_SIGNAL_X32_PLCWI", '1', STANDBY_SIGNAL_X32_PLCWI, test_failed);
  SEND_32_STANDBY_CTRL_WORDS_PLIF <= '0';
  wait for 10 us;
  --------------------------------------
  -- TEST 3:Loss Signal Control Word  --
  --------------------------------------
  -- test LOST_LIGNAL
  SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF      <= '1';
  LOST_CAUSE_MIB                          <= "11";
  wait until falling_edge(CLK);
  for i in 0 to 15 loop
    wait until falling_edge(CLK);
    check_equal("Test 3:Loss Signal Control Word : DATA_TX_PLCWI i="& integer'image(i)    ,    "000000" & "11" & C_LOST_SIG_WORD & "000000" & "11" & C_LOST_SIG_WORD, DATA_TX_PLCWI,        test_failed);
    check_equal("Test 3:Loss Signal Control Word : VALID_K_CHARAC_PLCWI i="& integer'image(i), x"11",                                                                   VALID_K_CHARAC_PLCWI, test_failed);
    check      ("Test 3:Loss Signal Control Word : NEW_DATA_PLCWI i="& integer'image(i),       '1' ,                                                                    NEW_DATA_PLCWI,       test_failed);
    check      ("Test 3:Loss Signal Control Word : LOST_SIGNAL_X32_PLCWI i="& integer'image(i),      '0' ,                                                                    LOST_SIGNAL_X32_PLCWI,      test_failed);
  end loop;
  wait until falling_edge(CLK);
  check      ("Test 3:Loss Signal Control Word : LOST_SIGNAL_X32_PLCWI", '1', LOST_SIGNAL_X32_PLCWI, test_failed);
  SEND_32_LOSS_SIGNAL_CTRL_WORDS_PLIF      <= '0';
  ------------------------------------------------------------
  --                       END TEST                         --
  ------------------------------------------------------------
  log_test_result(test_failed);

  wait;
end process;

end tb;