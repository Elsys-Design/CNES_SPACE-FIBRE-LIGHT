// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_PLLE4_ADV_DEFINES_VH
`else
`define B_PLLE4_ADV_DEFINES_VH

// Look-up table parameters
//

`define PLLE4_ADV_ADDR_N  24
`define PLLE4_ADV_ADDR_SZ 32
`define PLLE4_ADV_DATA_SZ 72

// Attribute addresses
//

`define PLLE4_ADV__CLKFBOUT_MULT    32'h00000000
`define PLLE4_ADV__CLKFBOUT_MULT_SZ 32

`define PLLE4_ADV__CLKFBOUT_PHASE    32'h00000001
`define PLLE4_ADV__CLKFBOUT_PHASE_SZ 64

`define PLLE4_ADV__CLKIN_FREQ_MAX    32'h00000002
`define PLLE4_ADV__CLKIN_FREQ_MAX_SZ 64

`define PLLE4_ADV__CLKIN_FREQ_MIN    32'h00000003
`define PLLE4_ADV__CLKIN_FREQ_MIN_SZ 64

`define PLLE4_ADV__CLKIN_PERIOD    32'h00000004
`define PLLE4_ADV__CLKIN_PERIOD_SZ 64

`define PLLE4_ADV__CLKOUT0_DIVIDE    32'h00000005
`define PLLE4_ADV__CLKOUT0_DIVIDE_SZ 32

`define PLLE4_ADV__CLKOUT0_DUTY_CYCLE    32'h00000006
`define PLLE4_ADV__CLKOUT0_DUTY_CYCLE_SZ 64

`define PLLE4_ADV__CLKOUT0_PHASE    32'h00000007
`define PLLE4_ADV__CLKOUT0_PHASE_SZ 64

`define PLLE4_ADV__CLKOUT1_DIVIDE    32'h00000008
`define PLLE4_ADV__CLKOUT1_DIVIDE_SZ 32

`define PLLE4_ADV__CLKOUT1_DUTY_CYCLE    32'h00000009
`define PLLE4_ADV__CLKOUT1_DUTY_CYCLE_SZ 64

`define PLLE4_ADV__CLKOUT1_PHASE    32'h0000000a
`define PLLE4_ADV__CLKOUT1_PHASE_SZ 64

`define PLLE4_ADV__CLKOUTPHY_MODE    32'h0000000b
`define PLLE4_ADV__CLKOUTPHY_MODE_SZ 64

`define PLLE4_ADV__CLKPFD_FREQ_MAX    32'h0000000c
`define PLLE4_ADV__CLKPFD_FREQ_MAX_SZ 64

`define PLLE4_ADV__CLKPFD_FREQ_MIN    32'h0000000d
`define PLLE4_ADV__CLKPFD_FREQ_MIN_SZ 64

`define PLLE4_ADV__COMPENSATION    32'h0000000e
`define PLLE4_ADV__COMPENSATION_SZ 72

`define PLLE4_ADV__DIVCLK_DIVIDE    32'h0000000f
`define PLLE4_ADV__DIVCLK_DIVIDE_SZ 32

`define PLLE4_ADV__IS_CLKFBIN_INVERTED    32'h00000010
`define PLLE4_ADV__IS_CLKFBIN_INVERTED_SZ 1

`define PLLE4_ADV__IS_CLKIN_INVERTED    32'h00000011
`define PLLE4_ADV__IS_CLKIN_INVERTED_SZ 1

`define PLLE4_ADV__IS_PWRDWN_INVERTED    32'h00000012
`define PLLE4_ADV__IS_PWRDWN_INVERTED_SZ 1

`define PLLE4_ADV__IS_RST_INVERTED    32'h00000013
`define PLLE4_ADV__IS_RST_INVERTED_SZ 1

`define PLLE4_ADV__REF_JITTER    32'h00000014
`define PLLE4_ADV__REF_JITTER_SZ 64

`define PLLE4_ADV__STARTUP_WAIT    32'h00000015
`define PLLE4_ADV__STARTUP_WAIT_SZ 40

`define PLLE4_ADV__VCOCLK_FREQ_MAX    32'h00000016
`define PLLE4_ADV__VCOCLK_FREQ_MAX_SZ 64

`define PLLE4_ADV__VCOCLK_FREQ_MIN    32'h00000017
`define PLLE4_ADV__VCOCLK_FREQ_MIN_SZ 64

`endif  // B_PLLE4_ADV_DEFINES_VH