// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_CPM5_DEFINES_VH
`else
`define B_CPM5_DEFINES_VH

// Look-up table parameters
//

`define CPM5_ADDR_N  21
`define CPM5_ADDR_SZ 32
`define CPM5_DATA_SZ 120

// Attribute addresses
//

`define CPM5__CLKDIV0    32'h00000000
`define CPM5__CLKDIV0_SZ 4

`define CPM5__CLKDIV1    32'h00000001
`define CPM5__CLKDIV1_SZ 4

`define CPM5__CPM5_DPLL0INT_DIVOUT    32'h00000002
`define CPM5__CPM5_DPLL0INT_DIVOUT_SZ 4

`define CPM5__CPM5_DPLL1INT_DIVOUT    32'h00000003
`define CPM5__CPM5_DPLL1INT_DIVOUT_SZ 4

`define CPM5__CPM5_MODE_0    32'h00000004
`define CPM5__CPM5_MODE_0_SZ 120

`define CPM5__CPM5_MODE_1    32'h00000005
`define CPM5__CPM5_MODE_1_SZ 120

`define CPM5__CXS0_MODE    32'h00000006
`define CPM5__CXS0_MODE_SZ 56

`define CPM5__CXS1_MODE    32'h00000007
`define CPM5__CXS1_MODE_SZ 56

`define CPM5__DPLL0_DESKEW_DELAY    32'h00000008
`define CPM5__DPLL0_DESKEW_DELAY_SZ 6

`define CPM5__DPLL0_DESKEW_DELAY_EN    32'h00000009
`define CPM5__DPLL0_DESKEW_DELAY_EN_SZ 40

`define CPM5__DPLL0_DESKEW_DELAY_PATH    32'h0000000a
`define CPM5__DPLL0_DESKEW_DELAY_PATH_SZ 40

`define CPM5__DPLL0_DESKEW_EN    32'h0000000b
`define CPM5__DPLL0_DESKEW_EN_SZ 40

`define CPM5__DPLL1_DESKEW_DELAY    32'h0000000c
`define CPM5__DPLL1_DESKEW_DELAY_SZ 6

`define CPM5__DPLL1_DESKEW_DELAY_EN    32'h0000000d
`define CPM5__DPLL1_DESKEW_DELAY_EN_SZ 40

`define CPM5__DPLL1_DESKEW_DELAY_PATH    32'h0000000e
`define CPM5__DPLL1_DESKEW_DELAY_PATH_SZ 40

`define CPM5__DPLL1_DESKEW_EN    32'h0000000f
`define CPM5__DPLL1_DESKEW_EN_SZ 40

`define CPM5__LINK_SPEED_0    32'h00000010
`define CPM5__LINK_SPEED_0_SZ 48

`define CPM5__LINK_SPEED_1    32'h00000011
`define CPM5__LINK_SPEED_1_SZ 48

`define CPM5__LINK_WIDTH_0    32'h00000012
`define CPM5__LINK_WIDTH_0_SZ 5

`define CPM5__LINK_WIDTH_1    32'h00000013
`define CPM5__LINK_WIDTH_1_SZ 4

`define CPM5__SIM_CPM_CDO_FILE_NAME    32'h00000014
`define CPM5__SIM_CPM_CDO_FILE_NAME_SZ 88

`endif  // B_CPM5_DEFINES_VH