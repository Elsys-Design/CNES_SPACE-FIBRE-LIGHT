-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 04/07/2025
--
-- Description : This is the testbench of the ppl_64_rx_sync_fsm module
----------------------------------------------------------------------------
LIBRARY ieee ;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

library work;
use work.pkg_simu.all;

entity tb_ppl_64_rx_sync_fsm is
end entity;

architecture tb of tb_ppl_64_rx_sync_fsm is
  component ppl_64_rx_sync_fsm is
    port(
      RST_N                            : in  std_logic;                                            --! global reset
      CLK                              : in  std_logic;                                            --! Clock generated by GTY IP
      -- FROM Data-link layer
      LANE_RESET_DL                    : in  std_logic;                                            --! Lane reset command from Data-Link Layer.
      -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
      DATA_RX_PLRSF                    : out std_logic_vector(C_DATA_LENGTH-1  downto 0);          --! 64-bit data to lane_ctrl_word_detect
      VALID_K_CHARAC_PLRSF             : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);  --! 8-bit valid K character flags to lane_ctrl_word_detect
      DATA_RDY_PLRSF                   : out std_logic;                                            --! Data valid flag to lane_ctrl_word_detect
      -- ppl_64_word_alignment (PLWA) interface
      DATA_RX_PLWA                     : in  std_logic_vector(C_DATA_LENGTH-1  downto 0);          --! 64-bit data from GTY IP
      VALID_K_CHARAC_PLWA              : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);  --! 8-bit valid K character flags from GTY IP
      INVALID_CHAR_PLWA                : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);  --! Invalid character flags from GTY IP
      DISPARITY_ERR_PLWA               : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);  --! Disparity error flags from GTY IP
      RX_WORD_IS_ALIGNED_PLWA          : in  std_logic;                                            --! RX word realign from GTY IP
      COMMA_DET_PLWA                   : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);  --! Flag indicates that a comma is detected on the word receive
      -- PARAMETERS (MIB)
      LANE_RESET                       : in  std_logic                                             --! Asserts or de-asserts LaneReset for the lane
    );
   end component;


---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
constant periode                        : time := 13.334 ns;

signal RST_N                            : std_logic := '0';
signal CLK                              : std_logic := '0';
-- FROM Data-link layer
signal LANE_RESET_DL                    : std_logic := '0';
-- TO lane_ctrl_word_detection
signal DATA_RX_PLRSF                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
signal VALID_K_CHARAC_PLRSF          : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0);
signal DATA_RDY_PLRSF                : std_logic;
-- FROM MANUFACTURER IP
signal DATA_RX_PLWA                  : std_logic_vector(C_DATA_LENGTH-1 downto 0)          := (others => '0');
signal VALID_K_CHARAC_PLWA           : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0) := (others => '0');
signal INVALID_CHAR_PLWA             : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0) := (others => '0');
signal DISPARITY_ERR_PLWA            : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0) := (others => '0');
signal RX_WORD_IS_ALIGNED_PLWA         : std_logic                                           := '1';
signal COMMA_DET_PLWA                : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1  downto 0) := (others => '0');
-- PARAMETERS
signal LANE_RESET                       : std_logic                                           := '0';

begin
----------------------------------------------------------------------------
-- Instantiation
----------------------------------------------------------------------------
DUT : ppl_64_rx_sync_fsm
   port map(
      RST_N                         => RST_N,
      CLK                           => CLK,
      -- FROM Data-link layer
      LANE_RESET_DL                 => LANE_RESET_DL,
      -- TO lane_ctrl_word_detection
      DATA_RX_PLRSF                 => DATA_RX_PLRSF,
      VALID_K_CHARAC_PLRSF          => VALID_K_CHARAC_PLRSF,
      DATA_RDY_PLRSF                => DATA_RDY_PLRSF,
      -- FROM MANUFACTURER IP
      DATA_RX_PLWA                  => DATA_RX_PLWA,
      VALID_K_CHARAC_PLWA           => VALID_K_CHARAC_PLWA,
      INVALID_CHAR_PLWA             => INVALID_CHAR_PLWA,
      DISPARITY_ERR_PLWA            => DISPARITY_ERR_PLWA,
      RX_WORD_IS_ALIGNED_PLWA       => RX_WORD_IS_ALIGNED_PLWA,
      COMMA_DET_PLWA                => COMMA_DET_PLWA,
      -- PARAMETERS
      LANE_RESET                    => LANE_RESET
      );


-- generate clock 75 MHz
horloge : process
begin
   CLK   <= not CLK;
   wait for periode/2;
end process;
----------------------------------------------------------------------------
-- Scenario
----------------------------------------------------------------------------
scenario : process
  variable test_failed : boolean := false;
begin

   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 20 us;
   ------------------------------------------------------------
   --   Test 0: Transition LOST_SYNC_ST                        --
   ------------------------------------------------------------
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   check_equal("Test 0: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 0: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 0: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 0: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 0: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 0: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   DATA_RX_PLWA         <= (others => '0');
   VALID_K_CHARAC_PLWA  <= (others => '0');
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 1: Transition LOST_SYNC_ST to CHECK_SYNC_ST       --
   ------------------------------------------------------------
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   check_equal("Test 1: DATA_RX_PLRSF_ERR"       , x"2222222211223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 1: VALID_K_CHARAC_PLRSF_ERR", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= (others => '0');
   VALID_K_CHARAC_PLWA  <= (others => '0');
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 2: LANE_RESET CHECK_SYNC_ST to LOST_SYNC_ST     --
   ------------------------------------------------------------
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   -- to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   --CHECK_SYNC_ST to LOST_SYNC_ST
   LANE_RESET  <= '1';
   wait until rising_edge(CLK);
   LANE_RESET  <= '0';
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   check_equal("Test 2: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 2: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 3: LANE_RESET READY_ST to LOST_SYNC_ST          --
   ------------------------------------------------------------
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   LANE_RESET  <= '1';
   wait until rising_edge(CLK);
   LANE_RESET  <= '0';
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   check_equal("Test 3: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 3: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= (others => '0');
   VALID_K_CHARAC_PLWA  <= (others => '0');
   wait for 10 us;
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 4 : LANE_RESET_DL CHECK_SYNC_ST to LOST_SYNC_ST    --
   ------------------------------------------------------------
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   LANE_RESET_DL  <= '1';
   wait until rising_edge(CLK);
   LANE_RESET_DL  <= '0';
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   check_equal("Test 4: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 4: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= (others => '0');
   VALID_K_CHARAC_PLWA  <= (others => '0');
   wait for 10 us;
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 5 : LANE_RESET_DL READY_ST to LOST_SYNC_ST      --
   ------------------------------------------------------------
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   LANE_RESET_DL  <= '1';
   wait until rising_edge(CLK);
   LANE_RESET_DL  <= '0';
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   check_equal("Test 5: DATA_RX_PLRSF_ERR"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 5: VALID_K_CHARAC_PLRSF_ERR", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= (others => '0');
   VALID_K_CHARAC_PLWA  <= (others => '0');
   wait for 10 us;
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 6: CHECK_SYNC_ST 1st word of the data bus wrong,  --
   --         only the second is valid => READY_ST           --
   ------------------------------------------------------------
   -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 10 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"01";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"0F";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"02";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_1"       , x"2222222200000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_1", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"0F";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"03";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_2"       , x"3333333300000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_2", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"0F";
   DATA_RX_PLWA         <= x"55555555DDEEFF00";
   VALID_K_CHARAC_PLWA  <= x"04";
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_3"       , x"4444444400000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_3", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"0F";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"6666666611223344";
   VALID_K_CHARAC_PLWA  <= x"05";
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_4"       , x"5555555500000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_4", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_5"       , x"6666666600000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_5", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 6: DATA_RX_PLRSF_ERR_5_6"       , x"6666666611223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 6: VALID_K_CHARAC_PLRSF_ERR_5_6", x"05",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 7: CHECK_SYNC_ST 2nd word of the data bus wrong,  --
   --         only the first one is valid => CHECK_SYNC_ST   --
   ------------------------------------------------------------
   -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 10 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"10";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"20";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_1"       , x"0000000011223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"F0";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"30";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_2"       , x"0000000055667788", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_2", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"55555555DDEEFF00";
   VALID_K_CHARAC_PLWA  <= x"40";
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_3"       , x"0000000099AABBCC", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_3", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"F0";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"6666666611223344";
   VALID_K_CHARAC_PLWA  <= x"05";
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_4"       , x"00000000DDEEFF00", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_4", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_5"       , x"0000000011223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_5", x"15",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 7: DATA_RX_PLRSF_ERR_5_6"       , x"6666666611223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 7: VALID_K_CHARAC_PLRSF_ERR_5_6", x"05",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 8: CHECK_SYNC_ST 2 words of the data bus wrong    --
   --         => LOST_SYNC_ST                                --
   ------------------------------------------------------------
   -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 10 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"11";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= x"01";
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_1"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"FF";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_2"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_2", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_3"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_3", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_4"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_4", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_5"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_5", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 8: DATA_RX_PLRSF_ERR_5_6"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 8: VALID_K_CHARAC_PLRSF_ERR_5_6", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 9 : READY_ST 1st word of the data bus wrong,     --
   --         only the second is valid => READY_ST           --
   ------------------------------------------------------------
      -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 9 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"01";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"0F";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"02";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_1"       , x"2222222200000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_1", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"0F";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"03";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_2"       , x"3333333300000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_2", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"0F";
   DATA_RX_PLWA         <= x"55555555DDEEFF00";
   VALID_K_CHARAC_PLWA  <= x"04";
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_3"       , x"4444444400000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_3", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"0F";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"6666666611223344";
   VALID_K_CHARAC_PLWA  <= x"05";
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_4"       , x"5555555500000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_4", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_5"       , x"6666666600000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_5", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 9: DATA_RX_PLRSF_ERR_5_6"       , x"6666666611223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 9: VALID_K_CHARAC_PLRSF_ERR_5_6", x"05",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 10 : READY_ST 2nd word of the data bus wrong,     --
   --         only the first one is valid => CHECK_SYNC_ST   --
   ------------------------------------------------------------
      -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 10 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"10";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"20";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_1"       , x"0000000011223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"F0";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"30";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_2"       , x"0000000055667788", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_2", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= (others => '0');
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"55555555DDEEFF00";
   VALID_K_CHARAC_PLWA  <= x"40";
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_3"       , x"0000000099AABBCC", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_3", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"F0";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"6666666611223344";
   VALID_K_CHARAC_PLWA  <= x"05";
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_4"       , x"00000000DDEEFF00", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_4", x"10",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_5"       , x"0000000011223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_5", x"15",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 10: DATA_RX_PLRSF_ERR_5_6"       , x"6666666611223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 10: VALID_K_CHARAC_PLRSF_ERR_5_6", x"05",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   -- Test 11 : READY_ST 2 words of the data bus wrong       --
   --         => LOST_SYNC_ST                                --
   ------------------------------------------------------------
      -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   wait until rising_edge(CLK);
   wait for 10 us;
   wait until rising_edge(CLK);     -- 1st word with error gen
   INVALID_CHAR_PLWA    <= x"11";
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 2nd word with errors gen
   INVALID_CHAR_PLWA    <= x"01";
   DISPARITY_ERR_PLWA   <= x"F0";
   DATA_RX_PLWA         <= x"3333333355667788";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 3rd word with errors gen and 1st word with error check
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_1"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA    <= x"FF";
   DISPARITY_ERR_PLWA   <= (others => '0');
   DATA_RX_PLWA         <= x"4444444499AABBCC";
   VALID_K_CHARAC_PLWA  <= x"00";
   wait until rising_edge(CLK);     -- 4nd word with errors gen and 2nd word with error check
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_2"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_2", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);     -- 5th word with errors gen and 3rd word with error check
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_3"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_3", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);-- 4th word with error check
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_4"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_4", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   INVALID_CHAR_PLWA  <= (others => '0');
   DISPARITY_ERR_PLWA <= (others => '0');
   wait until rising_edge(CLK);-- 5th word with error check
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_5"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_5", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 11: DATA_RX_PLRSF_ERR_5_6"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 11: VALID_K_CHARAC_PLRSF_ERR_5_6", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 12 : Realign CHECK_SYNC_ST to LOST_SYNC_ST      --
   ------------------------------------------------------------
   -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   check_equal("Test 12: DATA_RX_PLRSF_ERR_12_1"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 12: VALID_K_CHARAC_PLRSF_ERR_12_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
      -- CHECK_SYNC_ST to LOST_SYNC_ST
   RX_WORD_IS_ALIGNED_PLWA <= '0';
   wait until rising_edge(CLK);
   check_equal("Test 12: DATA_RX_PLRSF_ERR_12_2"       , x"2222222211223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 12: VALID_K_CHARAC_PLRSF_ERR_12_2", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 12: DATA_RX_PLRSF_ERR_12_3"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 12: VALID_K_CHARAC_PLRSF_ERR_12_3", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   -- Reset
   RX_WORD_IS_ALIGNED_PLWA <= '1';
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --   Test 13 : Realign READY_ST to LOST_SYNC_ST           --
   ------------------------------------------------------------
    -- LOST_SYNC_ST to CHECK_SYNC_ST
   COMMA_DET_PLWA <= "00000001";
   wait until rising_edge(CLK);
   COMMA_DET_PLWA <= (others => '0');
   check_equal("Test 13: DATA_RX_PLRSF_ERR_13_1"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 13: VALID_K_CHARAC_PLRSF_ERR_13_1", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= x"2222222211223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   wait until rising_edge(CLK);
   -- CHECK_SYNC_ST to READY_ST
   check_equal("Test 13: DATA_RX_PLRSF_ERR_13_2"       , x"2222222211223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 13: VALID_K_CHARAC_PLRSF_ERR_13_2", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   DATA_RX_PLWA         <= x"1111111111223344";
   VALID_K_CHARAC_PLWA  <= x"01";
   wait until rising_edge(CLK);
   -- READY_ST to LOST_SYNC_ST
   RX_WORD_IS_ALIGNED_PLWA <= '0';
   check_equal("Test 13: DATA_RX_PLRSF_ERR_13_3"       , x"2222222211223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 13: VALID_K_CHARAC_PLRSF_ERR_13_3", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 13: DATA_RX_PLRSF_ERR_13_4"       , x"1111111111223344", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 13: VALID_K_CHARAC_PLRSF_ERR_13_4", x"01",               VALID_K_CHARAC_PLRSF, test_failed);
   wait until rising_edge(CLK);
   check_equal("Test 13: DATA_RX_PLRSF_ERR_13_5"       , x"0000000000000000", DATA_RX_PLRSF,        test_failed);
   check_equal("Test 13: VALID_K_CHARAC_PLRSF_ERR_13_5", x"11",               VALID_K_CHARAC_PLRSF, test_failed);
   -- Reset
   wait for 10 us;
   RST_N <= '0';
   wait for 10 us;
   wait until rising_edge(CLK);
   RST_N <= '1';
   wait for 10 us;
   ------------------------------------------------------------
   --                       END TEST                         --
   ------------------------------------------------------------
   log_test_result(test_failed);


   wait;
end process;

end tb;