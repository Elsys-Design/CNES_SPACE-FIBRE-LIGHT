`include "B_CLOCK_MOD_IRI_IMR_defines.vh"

reg [`CLOCK_MOD_IRI_IMR_DATA_SZ-1:0] ATTR [0:`CLOCK_MOD_IRI_IMR_ADDR_N-1];
reg [`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_COE_SZ-1:0] CLK_DLY_VAL_COE_REG = CLK_DLY_VAL_COE;
reg [`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_IMUX_SZ-1:0] CLK_DLY_VAL_IMUX_REG = CLK_DLY_VAL_IMUX;
reg [`CLOCK_MOD_IRI_IMR__CLK_EN_SZ:1] CLK_EN_REG = CLK_EN;
reg [`CLOCK_MOD_IRI_IMR__IMUX_CLK1_SEL_SZ:1] IMUX_CLK1_SEL_REG = IMUX_CLK1_SEL;
reg [`CLOCK_MOD_IRI_IMR__IMUX_CLK2_SEL_SZ:1] IMUX_CLK2_SEL_REG = IMUX_CLK2_SEL;

initial begin
  ATTR[`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_COE] = CLK_DLY_VAL_COE;
  ATTR[`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_IMUX] = CLK_DLY_VAL_IMUX;
  ATTR[`CLOCK_MOD_IRI_IMR__CLK_EN] = CLK_EN;
  ATTR[`CLOCK_MOD_IRI_IMR__IMUX_CLK1_SEL] = IMUX_CLK1_SEL;
  ATTR[`CLOCK_MOD_IRI_IMR__IMUX_CLK2_SEL] = IMUX_CLK2_SEL;
end

always @(trig_attr) begin
  CLK_DLY_VAL_COE_REG = ATTR[`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_COE];
  CLK_DLY_VAL_IMUX_REG = ATTR[`CLOCK_MOD_IRI_IMR__CLK_DLY_VAL_IMUX];
  CLK_EN_REG = ATTR[`CLOCK_MOD_IRI_IMR__CLK_EN];
  IMUX_CLK1_SEL_REG = ATTR[`CLOCK_MOD_IRI_IMR__IMUX_CLK1_SEL];
  IMUX_CLK2_SEL_REG = ATTR[`CLOCK_MOD_IRI_IMR__IMUX_CLK2_SEL];
end

// procedures to override, read attribute values

task write_attr;
  input  [`CLOCK_MOD_IRI_IMR_ADDR_SZ-1:0] addr;
  input  [`CLOCK_MOD_IRI_IMR_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`CLOCK_MOD_IRI_IMR_DATA_SZ-1:0] read_attr;
  input  [`CLOCK_MOD_IRI_IMR_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
