// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSPCPLX_DEFINES_VH
`else
`define B_DSPCPLX_DEFINES_VH

// Look-up table parameters
//

`define DSPCPLX_ADDR_N  75
`define DSPCPLX_ADDR_SZ 32
`define DSPCPLX_DATA_SZ 120

// Attribute addresses
//

`define DSPCPLX__ACASCREG_IM    32'h00000000
`define DSPCPLX__ACASCREG_IM_SZ 32

`define DSPCPLX__ACASCREG_RE    32'h00000001
`define DSPCPLX__ACASCREG_RE_SZ 32

`define DSPCPLX__ADREG    32'h00000002
`define DSPCPLX__ADREG_SZ 32

`define DSPCPLX__ALUMODEREG_IM    32'h00000003
`define DSPCPLX__ALUMODEREG_IM_SZ 32

`define DSPCPLX__ALUMODEREG_RE    32'h00000004
`define DSPCPLX__ALUMODEREG_RE_SZ 32

`define DSPCPLX__AREG_IM    32'h00000005
`define DSPCPLX__AREG_IM_SZ 32

`define DSPCPLX__AREG_RE    32'h00000006
`define DSPCPLX__AREG_RE_SZ 32

`define DSPCPLX__AUTORESET_PATDET_IM    32'h00000007
`define DSPCPLX__AUTORESET_PATDET_IM_SZ 120

`define DSPCPLX__AUTORESET_PATDET_RE    32'h00000008
`define DSPCPLX__AUTORESET_PATDET_RE_SZ 120

`define DSPCPLX__AUTORESET_PRIORITY_IM    32'h00000009
`define DSPCPLX__AUTORESET_PRIORITY_IM_SZ 40

`define DSPCPLX__AUTORESET_PRIORITY_RE    32'h0000000a
`define DSPCPLX__AUTORESET_PRIORITY_RE_SZ 40

`define DSPCPLX__A_INPUT_IM    32'h0000000b
`define DSPCPLX__A_INPUT_IM_SZ 56

`define DSPCPLX__A_INPUT_RE    32'h0000000c
`define DSPCPLX__A_INPUT_RE_SZ 56

`define DSPCPLX__BCASCREG_IM    32'h0000000d
`define DSPCPLX__BCASCREG_IM_SZ 32

`define DSPCPLX__BCASCREG_RE    32'h0000000e
`define DSPCPLX__BCASCREG_RE_SZ 32

`define DSPCPLX__BREG_IM    32'h0000000f
`define DSPCPLX__BREG_IM_SZ 32

`define DSPCPLX__BREG_RE    32'h00000010
`define DSPCPLX__BREG_RE_SZ 32

`define DSPCPLX__B_INPUT_IM    32'h00000011
`define DSPCPLX__B_INPUT_IM_SZ 56

`define DSPCPLX__B_INPUT_RE    32'h00000012
`define DSPCPLX__B_INPUT_RE_SZ 56

`define DSPCPLX__CARRYINREG_IM    32'h00000013
`define DSPCPLX__CARRYINREG_IM_SZ 32

`define DSPCPLX__CARRYINREG_RE    32'h00000014
`define DSPCPLX__CARRYINREG_RE_SZ 32

`define DSPCPLX__CARRYINSELREG_IM    32'h00000015
`define DSPCPLX__CARRYINSELREG_IM_SZ 32

`define DSPCPLX__CARRYINSELREG_RE    32'h00000016
`define DSPCPLX__CARRYINSELREG_RE_SZ 32

`define DSPCPLX__CONJUGATEREG_A    32'h00000017
`define DSPCPLX__CONJUGATEREG_A_SZ 32

`define DSPCPLX__CONJUGATEREG_B    32'h00000018
`define DSPCPLX__CONJUGATEREG_B_SZ 32

`define DSPCPLX__CREG_IM    32'h00000019
`define DSPCPLX__CREG_IM_SZ 32

`define DSPCPLX__CREG_RE    32'h0000001a
`define DSPCPLX__CREG_RE_SZ 32

`define DSPCPLX__IS_ALUMODE_IM_INVERTED    32'h0000001b
`define DSPCPLX__IS_ALUMODE_IM_INVERTED_SZ 4

`define DSPCPLX__IS_ALUMODE_RE_INVERTED    32'h0000001c
`define DSPCPLX__IS_ALUMODE_RE_INVERTED_SZ 4

`define DSPCPLX__IS_ASYNC_RST_INVERTED    32'h0000001d
`define DSPCPLX__IS_ASYNC_RST_INVERTED_SZ 1

`define DSPCPLX__IS_CARRYIN_IM_INVERTED    32'h0000001e
`define DSPCPLX__IS_CARRYIN_IM_INVERTED_SZ 1

`define DSPCPLX__IS_CARRYIN_RE_INVERTED    32'h0000001f
`define DSPCPLX__IS_CARRYIN_RE_INVERTED_SZ 1

`define DSPCPLX__IS_CLK_INVERTED    32'h00000020
`define DSPCPLX__IS_CLK_INVERTED_SZ 1

`define DSPCPLX__IS_CONJUGATE_A_INVERTED    32'h00000021
`define DSPCPLX__IS_CONJUGATE_A_INVERTED_SZ 1

`define DSPCPLX__IS_CONJUGATE_B_INVERTED    32'h00000022
`define DSPCPLX__IS_CONJUGATE_B_INVERTED_SZ 1

`define DSPCPLX__IS_OPMODE_IM_INVERTED    32'h00000023
`define DSPCPLX__IS_OPMODE_IM_INVERTED_SZ 9

`define DSPCPLX__IS_OPMODE_RE_INVERTED    32'h00000024
`define DSPCPLX__IS_OPMODE_RE_INVERTED_SZ 9

`define DSPCPLX__IS_RSTAD_INVERTED    32'h00000025
`define DSPCPLX__IS_RSTAD_INVERTED_SZ 1

`define DSPCPLX__IS_RSTALLCARRYIN_IM_INVERTED    32'h00000026
`define DSPCPLX__IS_RSTALLCARRYIN_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTALLCARRYIN_RE_INVERTED    32'h00000027
`define DSPCPLX__IS_RSTALLCARRYIN_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTALUMODE_IM_INVERTED    32'h00000028
`define DSPCPLX__IS_RSTALUMODE_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTALUMODE_RE_INVERTED    32'h00000029
`define DSPCPLX__IS_RSTALUMODE_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTA_IM_INVERTED    32'h0000002a
`define DSPCPLX__IS_RSTA_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTA_RE_INVERTED    32'h0000002b
`define DSPCPLX__IS_RSTA_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTB_IM_INVERTED    32'h0000002c
`define DSPCPLX__IS_RSTB_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTB_RE_INVERTED    32'h0000002d
`define DSPCPLX__IS_RSTB_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTCONJUGATE_A_INVERTED    32'h0000002e
`define DSPCPLX__IS_RSTCONJUGATE_A_INVERTED_SZ 1

`define DSPCPLX__IS_RSTCONJUGATE_B_INVERTED    32'h0000002f
`define DSPCPLX__IS_RSTCONJUGATE_B_INVERTED_SZ 1

`define DSPCPLX__IS_RSTCTRL_IM_INVERTED    32'h00000030
`define DSPCPLX__IS_RSTCTRL_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTCTRL_RE_INVERTED    32'h00000031
`define DSPCPLX__IS_RSTCTRL_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTC_IM_INVERTED    32'h00000032
`define DSPCPLX__IS_RSTC_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTC_RE_INVERTED    32'h00000033
`define DSPCPLX__IS_RSTC_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTM_IM_INVERTED    32'h00000034
`define DSPCPLX__IS_RSTM_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTM_RE_INVERTED    32'h00000035
`define DSPCPLX__IS_RSTM_RE_INVERTED_SZ 1

`define DSPCPLX__IS_RSTP_IM_INVERTED    32'h00000036
`define DSPCPLX__IS_RSTP_IM_INVERTED_SZ 1

`define DSPCPLX__IS_RSTP_RE_INVERTED    32'h00000037
`define DSPCPLX__IS_RSTP_RE_INVERTED_SZ 1

`define DSPCPLX__MASK_IM    32'h00000038
`define DSPCPLX__MASK_IM_SZ 58

`define DSPCPLX__MASK_RE    32'h00000039
`define DSPCPLX__MASK_RE_SZ 58

`define DSPCPLX__MREG_IM    32'h0000003a
`define DSPCPLX__MREG_IM_SZ 32

`define DSPCPLX__MREG_RE    32'h0000003b
`define DSPCPLX__MREG_RE_SZ 32

`define DSPCPLX__OPMODEREG_IM    32'h0000003c
`define DSPCPLX__OPMODEREG_IM_SZ 32

`define DSPCPLX__OPMODEREG_RE    32'h0000003d
`define DSPCPLX__OPMODEREG_RE_SZ 32

`define DSPCPLX__PATTERN_IM    32'h0000003e
`define DSPCPLX__PATTERN_IM_SZ 58

`define DSPCPLX__PATTERN_RE    32'h0000003f
`define DSPCPLX__PATTERN_RE_SZ 58

`define DSPCPLX__PREG_IM    32'h00000040
`define DSPCPLX__PREG_IM_SZ 32

`define DSPCPLX__PREG_RE    32'h00000041
`define DSPCPLX__PREG_RE_SZ 32

`define DSPCPLX__RESET_MODE    32'h00000042
`define DSPCPLX__RESET_MODE_SZ 40

`define DSPCPLX__RND_IM    32'h00000043
`define DSPCPLX__RND_IM_SZ 58

`define DSPCPLX__RND_RE    32'h00000044
`define DSPCPLX__RND_RE_SZ 58

`define DSPCPLX__SEL_MASK_IM    32'h00000045
`define DSPCPLX__SEL_MASK_IM_SZ 112

`define DSPCPLX__SEL_MASK_RE    32'h00000046
`define DSPCPLX__SEL_MASK_RE_SZ 112

`define DSPCPLX__SEL_PATTERN_IM    32'h00000047
`define DSPCPLX__SEL_PATTERN_IM_SZ 56

`define DSPCPLX__SEL_PATTERN_RE    32'h00000048
`define DSPCPLX__SEL_PATTERN_RE_SZ 56

`define DSPCPLX__USE_PATTERN_DETECT_IM    32'h00000049
`define DSPCPLX__USE_PATTERN_DETECT_IM_SZ 72

`define DSPCPLX__USE_PATTERN_DETECT_RE    32'h0000004a
`define DSPCPLX__USE_PATTERN_DETECT_RE_SZ 72

`endif  // B_DSPCPLX_DEFINES_VH