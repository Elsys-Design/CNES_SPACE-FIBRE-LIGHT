// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_BITSLICE_CONTROL_DEFINES_VH
`else
`define B_BITSLICE_CONTROL_DEFINES_VH

// Look-up table parameters
//

`define BITSLICE_CONTROL_ADDR_N  24
`define BITSLICE_CONTROL_ADDR_SZ 32
`define BITSLICE_CONTROL_DATA_SZ 152

// Attribute addresses
//

`define BITSLICE_CONTROL__CTRL_CLK    32'h00000000
`define BITSLICE_CONTROL__CTRL_CLK_SZ 64

`define BITSLICE_CONTROL__DIV_MODE    32'h00000001
`define BITSLICE_CONTROL__DIV_MODE_SZ 32

`define BITSLICE_CONTROL__EN_CLK_TO_EXT_NORTH    32'h00000002
`define BITSLICE_CONTROL__EN_CLK_TO_EXT_NORTH_SZ 56

`define BITSLICE_CONTROL__EN_CLK_TO_EXT_SOUTH    32'h00000003
`define BITSLICE_CONTROL__EN_CLK_TO_EXT_SOUTH_SZ 56

`define BITSLICE_CONTROL__EN_DYN_ODLY_MODE    32'h00000004
`define BITSLICE_CONTROL__EN_DYN_ODLY_MODE_SZ 40

`define BITSLICE_CONTROL__EN_OTHER_NCLK    32'h00000005
`define BITSLICE_CONTROL__EN_OTHER_NCLK_SZ 40

`define BITSLICE_CONTROL__EN_OTHER_PCLK    32'h00000006
`define BITSLICE_CONTROL__EN_OTHER_PCLK_SZ 40

`define BITSLICE_CONTROL__IDLY_VT_TRACK    32'h00000007
`define BITSLICE_CONTROL__IDLY_VT_TRACK_SZ 40

`define BITSLICE_CONTROL__INV_RXCLK    32'h00000008
`define BITSLICE_CONTROL__INV_RXCLK_SZ 40

`define BITSLICE_CONTROL__ODLY_VT_TRACK    32'h00000009
`define BITSLICE_CONTROL__ODLY_VT_TRACK_SZ 40

`define BITSLICE_CONTROL__QDLY_VT_TRACK    32'h0000000a
`define BITSLICE_CONTROL__QDLY_VT_TRACK_SZ 40

`define BITSLICE_CONTROL__READ_IDLE_COUNT    32'h0000000b
`define BITSLICE_CONTROL__READ_IDLE_COUNT_SZ 6

`define BITSLICE_CONTROL__REFCLK_SRC    32'h0000000c
`define BITSLICE_CONTROL__REFCLK_SRC_SZ 48

`define BITSLICE_CONTROL__ROUNDING_FACTOR    32'h0000000d
`define BITSLICE_CONTROL__ROUNDING_FACTOR_SZ 8

`define BITSLICE_CONTROL__RXGATE_EXTEND    32'h0000000e
`define BITSLICE_CONTROL__RXGATE_EXTEND_SZ 40

`define BITSLICE_CONTROL__RX_CLK_PHASE_N    32'h0000000f
`define BITSLICE_CONTROL__RX_CLK_PHASE_N_SZ 64

`define BITSLICE_CONTROL__RX_CLK_PHASE_P    32'h00000010
`define BITSLICE_CONTROL__RX_CLK_PHASE_P_SZ 64

`define BITSLICE_CONTROL__RX_GATING    32'h00000011
`define BITSLICE_CONTROL__RX_GATING_SZ 56

`define BITSLICE_CONTROL__SELF_CALIBRATE    32'h00000012
`define BITSLICE_CONTROL__SELF_CALIBRATE_SZ 56

`define BITSLICE_CONTROL__SERIAL_MODE    32'h00000013
`define BITSLICE_CONTROL__SERIAL_MODE_SZ 40

`define BITSLICE_CONTROL__SIM_DEVICE    32'h00000014
`define BITSLICE_CONTROL__SIM_DEVICE_SZ 152

`define BITSLICE_CONTROL__SIM_SPEEDUP    32'h00000015
`define BITSLICE_CONTROL__SIM_SPEEDUP_SZ 32

`define BITSLICE_CONTROL__SIM_VERSION    32'h00000016
`define BITSLICE_CONTROL__SIM_VERSION_SZ 64

`define BITSLICE_CONTROL__TX_GATING    32'h00000017
`define BITSLICE_CONTROL__TX_GATING_SZ 56

`endif  // B_BITSLICE_CONTROL_DEFINES_VH