----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module checks the validity of the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_desencapsulation is
  generic (
    G_VC_NUM       : integer := 8                                                  --! Number of virtual channel
 );
  port (
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- DBUFI interface
    DATA_DBUFI             : in std_logic_vector(C_DATA_LENGTH+C_BYTE_BY_WORD_LENGTH-1 downto 0);    -- Data read bus
    DATA_EN_DBUFI          : out  std_logic;                                -- Read command
    DATA_VLD_DBUFI         : in std_logic;                                -- Data valid
    -- DOBUF interface
    FCT_FAR_END_DDES       : out  std_logic_vector(G_VC_NUM-1 downto 0);    -- Data write bus
    MULT_DDES              : out  vc_mult_array(G_VC_NUM-1 downto 0);    -- Data write bus
    -- DIBUF interface
    DATA_DDES              : out  vc_data_k_array(G_VC_NUM downto 0);    -- Data & k write vc & broadcast
    DATA_EN_DDES           : out  std_logic_vector(G_VC_NUM downto 0);   -- Write command vc & broadcast
  );
end data_seq_check;

architecture rtl of data_desencapsulation is
---------------------------------------------------------
-----                  Declaration signals          -----
---------------------------------------------------------
signal data_in    : std_logic_vector(C_DATA_LENGTH+C_BYTE_BY_WORD_LENGTH-1 downto 0);
signal k_char_in  : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);

begin

  data_in   <= DATA_DBUFI(C_DATA_LENGTH-1 downto 0);
  k_char_in <= DATA_DBUFI(C_DATA_LENGTH+C_BYTE_BY_WORD_LENGTH-1 downto C_DATA_LENGTH);
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_seq_num
-- Description: Check the SEQ_NUM for each frame 
---------------------------------------------------------


end architecture rtl;