`include "B_HBM_SNGLBLI_INTF_AXI_TEST_defines.vh"

reg [`HBM_SNGLBLI_INTF_AXI_TEST_DATA_SZ-1:0] ATTR [0:`HBM_SNGLBLI_INTF_AXI_TEST_ADDR_N-1];
reg [40:1] APB_BYPASS_EN_REG = APB_BYPASS_EN;
reg [40:1] AXI_BYPASS_EN_REG = AXI_BYPASS_EN;
reg [40:1] CLK_SEL_REG = CLK_SEL;
reg [51:0] DBG_BYPASS_VAL_REG = DBG_BYPASS_VAL;
reg [40:1] DEBUG_MODE_REG = DEBUG_MODE;
reg [31:0] DFI_BYPASS_VAL_REG = DFI_BYPASS_VAL;
reg [40:1] MC_ENABLE_REG = MC_ENABLE;
reg [40:1] PHY_ENABLE_REG = PHY_ENABLE;
reg [40:1] SWITCH_ENABLE_REG = SWITCH_ENABLE;

initial begin
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__APB_BYPASS_EN] = APB_BYPASS_EN;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__AXI_BYPASS_EN] = AXI_BYPASS_EN;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__CLK_SEL] = CLK_SEL;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DBG_BYPASS_VAL] = DBG_BYPASS_VAL;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DEBUG_MODE] = DEBUG_MODE;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DFI_BYPASS_VAL] = DFI_BYPASS_VAL;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__MC_ENABLE] = MC_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__PHY_ENABLE] = PHY_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__SWITCH_ENABLE] = SWITCH_ENABLE;
end

always @(trig_attr) begin
  APB_BYPASS_EN_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__APB_BYPASS_EN];
  AXI_BYPASS_EN_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__AXI_BYPASS_EN];
  CLK_SEL_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__CLK_SEL];
  DBG_BYPASS_VAL_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DBG_BYPASS_VAL];
  DEBUG_MODE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DEBUG_MODE];
  DFI_BYPASS_VAL_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__DFI_BYPASS_VAL];
  MC_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__MC_ENABLE];
  PHY_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__PHY_ENABLE];
  SWITCH_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_AXI_TEST__SWITCH_ENABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`HBM_SNGLBLI_INTF_AXI_TEST_ADDR_SZ-1:0] addr;
  input  [`HBM_SNGLBLI_INTF_AXI_TEST_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`HBM_SNGLBLI_INTF_AXI_TEST_DATA_SZ-1:0] read_attr;
  input  [`HBM_SNGLBLI_INTF_AXI_TEST_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
