// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IBUF_INTERMDISABLE_DEFINES_VH
`else
`define B_IBUF_INTERMDISABLE_DEFINES_VH

// Look-up table parameters
//

`define IBUF_INTERMDISABLE_ADDR_N  4
`define IBUF_INTERMDISABLE_ADDR_SZ 32
`define IBUF_INTERMDISABLE_DATA_SZ 88

// Attribute addresses
//

`define IBUF_INTERMDISABLE__IBUF_LOW_PWR    32'h00000000
`define IBUF_INTERMDISABLE__IBUF_LOW_PWR_SZ 40

`define IBUF_INTERMDISABLE__IOSTANDARD    32'h00000001
`define IBUF_INTERMDISABLE__IOSTANDARD_SZ 56

`define IBUF_INTERMDISABLE__SIM_DEVICE    32'h00000002
`define IBUF_INTERMDISABLE__SIM_DEVICE_SZ 88

`define IBUF_INTERMDISABLE__USE_IBUFDISABLE    32'h00000003
`define IBUF_INTERMDISABLE__USE_IBUFDISABLE_SZ 40

`endif  // B_IBUF_INTERMDISABLE_DEFINES_VH