-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/03/2025
--
-- Description : This module computes the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

entity data_seq_compute is
port (
	CLK                   : in  std_logic;                                           --! Clock generated by GTY IP
  -- data_link_reset (DLRE) interface
  LINK_RESET_DLRE       : in  std_logic;                                           --! Link Reset command
  -- phy_plus_lane (PPL) interface
  LANE_ACTIVE_PPL       : in  std_logic;                                           --! Lane Active flag for the DATA Link Layer
	-- data_encapsulation (DENC) interface
	NEW_WORD_DENC         : in  std_logic;                                           --! New word flag associated with DATA_DENC
	DATA_DENC             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel from data_encapsulation
	VALID_K_CHARAC_DENC   : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K charachter valid in the 32-bit DATA_DENC vector
	TYPE_FRAME_DENC       : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Type of the frame associated with DATA_DENC
	END_FRAME_DENC        : in  std_logic;                                           --! End frame/control word associated with DATA_DENC
	SEQ_NUM_ACK_DENC      : in  std_logic_vector(7 downto 0);                        --! SEQ_NUM ACK value
	TRANS_POL_FLG_DENC    : in  std_logic;                                           --! Transmission polarity flag
	-- data_crc_compute (DCCHECK) interface
	NEW_WORD_DSCOM        : out std_logic;                                           --! New word flag associated with DATA_DSCOM
	DATA_DSCOM            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel to data_encapsulation
	VALID_K_CHARAC_DSCOM  : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K charachter valid in the 32-bit DATA_DSCOM vector
	TYPE_FRAME_DSCOM      : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Type of the frame associated with DATA_DSCOM
	END_FRAME_DSCOM       : out std_logic;                                           --! End frame/control word associated with DATA_DSCOM
	-- MIB interface
	SEQ_NUM_DSCOM         : out std_logic_vector(7 downto 0)                         --! Current SEQ_NUM value
  );
end data_seq_compute;

architecture rtl of data_seq_compute is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------

signal trans_seq_cnt    : unsigned(6 downto 0);
begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_seq_num_comp
-- Description: Computes the SEQ_NUM for each frame
---------------------------------------------------------
p_seq_num_comp: process(CLK)
begin
	if rising_edge(CLK)  then
    if LINK_RESET_DLRE ='1' then
	  	trans_seq_cnt        <= (others => '0'); -- Reset seq_num_cnt	on link reset
			NEW_WORD_DSCOM       <= '0';
			VALID_K_CHARAC_DSCOM <= (others => '0');
			TYPE_FRAME_DSCOM     <= (others => '0');
			END_FRAME_DSCOM      <= '0';
			DATA_DSCOM           <= (others => '0');
			SEQ_NUM_DSCOM        <= (others => '0');
		elsif LANE_ACTIVE_PPL= '1' then
			NEW_WORD_DSCOM       <= NEW_WORD_DENC;
			VALID_K_CHARAC_DSCOM <= VALID_K_CHARAC_DENC;
			TYPE_FRAME_DSCOM     <= TYPE_FRAME_DENC;
			END_FRAME_DSCOM      <= END_FRAME_DENC;
			if END_FRAME_DENC = '1' then -- control word or EDF or EBF
				if TYPE_FRAME_DENC = C_DATA_FRM then
					DATA_DSCOM      <= C_RESERVED_SYMB & C_RESERVED_SYMB & TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt+1) & DATA_DENC(7 downto 0);
					SEQ_NUM_DSCOM   <= TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt+1);
					trans_seq_cnt   <= trans_seq_cnt +1;
				elsif TYPE_FRAME_DENC = C_BC_FRM or TYPE_FRAME_DENC = C_FCT_FRM then
					DATA_DSCOM      <= C_RESERVED_SYMB & TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt+1) & DATA_DENC(15 downto 0);
					SEQ_NUM_DSCOM   <= TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt+1);
					trans_seq_cnt   <= trans_seq_cnt +1;
				elsif TYPE_FRAME_DENC = C_ACK_FRM or TYPE_FRAME_DENC = C_NACK_FRM then
					DATA_DSCOM      <= C_RESERVED_SYMB & SEQ_NUM_ACK_DENC & DATA_DENC(15 downto 0);
				else
					DATA_DSCOM      <= C_RESERVED_SYMB & TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt) & DATA_DENC(15 downto 0);
					SEQ_NUM_DSCOM   <= TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt);
				end if;
			elsif DATA_DENC(15 downto 0) = C_SIF_WORD and VALID_K_CHARAC_DENC(0)= '1' then -- SIF
				DATA_DSCOM      <= C_RESERVED_SYMB & TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt) & DATA_DENC(15 downto 0);
				SEQ_NUM_DSCOM   <= TRANS_POL_FLG_DENC & std_logic_vector(trans_seq_cnt);
			else
  	    DATA_DSCOM      <= DATA_DENC;
			end if;
		end if;
	end if;
end process p_seq_num_comp;

end architecture rtl;