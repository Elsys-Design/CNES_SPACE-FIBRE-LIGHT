// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_FPM_PIPEREG_DEFINES_VH
`else
`define B_DSP_FPM_PIPEREG_DEFINES_VH

// Look-up table parameters
//

`define DSP_FPM_PIPEREG_ADDR_N  6
`define DSP_FPM_PIPEREG_ADDR_SZ 32
`define DSP_FPM_PIPEREG_DATA_SZ 64

// Attribute addresses
//

`define DSP_FPM_PIPEREG__A_FPTYPE    32'h00000000
`define DSP_FPM_PIPEREG__A_FPTYPE_SZ 24

`define DSP_FPM_PIPEREG__B_D_FPTYPE    32'h00000001
`define DSP_FPM_PIPEREG__B_D_FPTYPE_SZ 24

`define DSP_FPM_PIPEREG__FPMPIPEREG    32'h00000002
`define DSP_FPM_PIPEREG__FPMPIPEREG_SZ 32

`define DSP_FPM_PIPEREG__IS_RSTFPMPIPE_INVERTED    32'h00000003
`define DSP_FPM_PIPEREG__IS_RSTFPMPIPE_INVERTED_SZ 1

`define DSP_FPM_PIPEREG__RESET_MODE    32'h00000004
`define DSP_FPM_PIPEREG__RESET_MODE_SZ 40

`define DSP_FPM_PIPEREG__USE_MULT    32'h00000005
`define DSP_FPM_PIPEREG__USE_MULT_SZ 64

`endif  // B_DSP_FPM_PIPEREG_DEFINES_VH