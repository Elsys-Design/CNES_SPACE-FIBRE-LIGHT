// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_RAMB36E2_DEFINES_VH
`else
`define B_RAMB36E2_DEFINES_VH

// Look-up table parameters
//

`define RAMB36E2_ADDR_N  179
`define RAMB36E2_ADDR_SZ 32
`define RAMB36E2_DATA_SZ 256

// Attribute addresses
//

`define RAMB36E2__CASCADE_ORDER_A    32'h00000000
`define RAMB36E2__CASCADE_ORDER_A_SZ 48

`define RAMB36E2__CASCADE_ORDER_B    32'h00000001
`define RAMB36E2__CASCADE_ORDER_B_SZ 48

`define RAMB36E2__CLOCK_DOMAINS    32'h00000002
`define RAMB36E2__CLOCK_DOMAINS_SZ 88

`define RAMB36E2__DOA_REG    32'h00000003
`define RAMB36E2__DOA_REG_SZ 32

`define RAMB36E2__DOB_REG    32'h00000004
`define RAMB36E2__DOB_REG_SZ 32

`define RAMB36E2__ENADDRENA    32'h00000005
`define RAMB36E2__ENADDRENA_SZ 40

`define RAMB36E2__ENADDRENB    32'h00000006
`define RAMB36E2__ENADDRENB_SZ 40

`define RAMB36E2__EN_ECC_PIPE    32'h00000007
`define RAMB36E2__EN_ECC_PIPE_SZ 40

`define RAMB36E2__EN_ECC_READ    32'h00000008
`define RAMB36E2__EN_ECC_READ_SZ 40

`define RAMB36E2__EN_ECC_WRITE    32'h00000009
`define RAMB36E2__EN_ECC_WRITE_SZ 40

`define RAMB36E2__INITP_00    32'h0000000a
`define RAMB36E2__INITP_00_SZ 256

`define RAMB36E2__INITP_01    32'h0000000b
`define RAMB36E2__INITP_01_SZ 256

`define RAMB36E2__INITP_02    32'h0000000c
`define RAMB36E2__INITP_02_SZ 256

`define RAMB36E2__INITP_03    32'h0000000d
`define RAMB36E2__INITP_03_SZ 256

`define RAMB36E2__INITP_04    32'h0000000e
`define RAMB36E2__INITP_04_SZ 256

`define RAMB36E2__INITP_05    32'h0000000f
`define RAMB36E2__INITP_05_SZ 256

`define RAMB36E2__INITP_06    32'h00000010
`define RAMB36E2__INITP_06_SZ 256

`define RAMB36E2__INITP_07    32'h00000011
`define RAMB36E2__INITP_07_SZ 256

`define RAMB36E2__INITP_08    32'h00000012
`define RAMB36E2__INITP_08_SZ 256

`define RAMB36E2__INITP_09    32'h00000013
`define RAMB36E2__INITP_09_SZ 256

`define RAMB36E2__INITP_0A    32'h00000014
`define RAMB36E2__INITP_0A_SZ 256

`define RAMB36E2__INITP_0B    32'h00000015
`define RAMB36E2__INITP_0B_SZ 256

`define RAMB36E2__INITP_0C    32'h00000016
`define RAMB36E2__INITP_0C_SZ 256

`define RAMB36E2__INITP_0D    32'h00000017
`define RAMB36E2__INITP_0D_SZ 256

`define RAMB36E2__INITP_0E    32'h00000018
`define RAMB36E2__INITP_0E_SZ 256

`define RAMB36E2__INITP_0F    32'h00000019
`define RAMB36E2__INITP_0F_SZ 256

`define RAMB36E2__INIT_00    32'h0000001a
`define RAMB36E2__INIT_00_SZ 256

`define RAMB36E2__INIT_01    32'h0000001b
`define RAMB36E2__INIT_01_SZ 256

`define RAMB36E2__INIT_02    32'h0000001c
`define RAMB36E2__INIT_02_SZ 256

`define RAMB36E2__INIT_03    32'h0000001d
`define RAMB36E2__INIT_03_SZ 256

`define RAMB36E2__INIT_04    32'h0000001e
`define RAMB36E2__INIT_04_SZ 256

`define RAMB36E2__INIT_05    32'h0000001f
`define RAMB36E2__INIT_05_SZ 256

`define RAMB36E2__INIT_06    32'h00000020
`define RAMB36E2__INIT_06_SZ 256

`define RAMB36E2__INIT_07    32'h00000021
`define RAMB36E2__INIT_07_SZ 256

`define RAMB36E2__INIT_08    32'h00000022
`define RAMB36E2__INIT_08_SZ 256

`define RAMB36E2__INIT_09    32'h00000023
`define RAMB36E2__INIT_09_SZ 256

`define RAMB36E2__INIT_0A    32'h00000024
`define RAMB36E2__INIT_0A_SZ 256

`define RAMB36E2__INIT_0B    32'h00000025
`define RAMB36E2__INIT_0B_SZ 256

`define RAMB36E2__INIT_0C    32'h00000026
`define RAMB36E2__INIT_0C_SZ 256

`define RAMB36E2__INIT_0D    32'h00000027
`define RAMB36E2__INIT_0D_SZ 256

`define RAMB36E2__INIT_0E    32'h00000028
`define RAMB36E2__INIT_0E_SZ 256

`define RAMB36E2__INIT_0F    32'h00000029
`define RAMB36E2__INIT_0F_SZ 256

`define RAMB36E2__INIT_10    32'h0000002a
`define RAMB36E2__INIT_10_SZ 256

`define RAMB36E2__INIT_11    32'h0000002b
`define RAMB36E2__INIT_11_SZ 256

`define RAMB36E2__INIT_12    32'h0000002c
`define RAMB36E2__INIT_12_SZ 256

`define RAMB36E2__INIT_13    32'h0000002d
`define RAMB36E2__INIT_13_SZ 256

`define RAMB36E2__INIT_14    32'h0000002e
`define RAMB36E2__INIT_14_SZ 256

`define RAMB36E2__INIT_15    32'h0000002f
`define RAMB36E2__INIT_15_SZ 256

`define RAMB36E2__INIT_16    32'h00000030
`define RAMB36E2__INIT_16_SZ 256

`define RAMB36E2__INIT_17    32'h00000031
`define RAMB36E2__INIT_17_SZ 256

`define RAMB36E2__INIT_18    32'h00000032
`define RAMB36E2__INIT_18_SZ 256

`define RAMB36E2__INIT_19    32'h00000033
`define RAMB36E2__INIT_19_SZ 256

`define RAMB36E2__INIT_1A    32'h00000034
`define RAMB36E2__INIT_1A_SZ 256

`define RAMB36E2__INIT_1B    32'h00000035
`define RAMB36E2__INIT_1B_SZ 256

`define RAMB36E2__INIT_1C    32'h00000036
`define RAMB36E2__INIT_1C_SZ 256

`define RAMB36E2__INIT_1D    32'h00000037
`define RAMB36E2__INIT_1D_SZ 256

`define RAMB36E2__INIT_1E    32'h00000038
`define RAMB36E2__INIT_1E_SZ 256

`define RAMB36E2__INIT_1F    32'h00000039
`define RAMB36E2__INIT_1F_SZ 256

`define RAMB36E2__INIT_20    32'h0000003a
`define RAMB36E2__INIT_20_SZ 256

`define RAMB36E2__INIT_21    32'h0000003b
`define RAMB36E2__INIT_21_SZ 256

`define RAMB36E2__INIT_22    32'h0000003c
`define RAMB36E2__INIT_22_SZ 256

`define RAMB36E2__INIT_23    32'h0000003d
`define RAMB36E2__INIT_23_SZ 256

`define RAMB36E2__INIT_24    32'h0000003e
`define RAMB36E2__INIT_24_SZ 256

`define RAMB36E2__INIT_25    32'h0000003f
`define RAMB36E2__INIT_25_SZ 256

`define RAMB36E2__INIT_26    32'h00000040
`define RAMB36E2__INIT_26_SZ 256

`define RAMB36E2__INIT_27    32'h00000041
`define RAMB36E2__INIT_27_SZ 256

`define RAMB36E2__INIT_28    32'h00000042
`define RAMB36E2__INIT_28_SZ 256

`define RAMB36E2__INIT_29    32'h00000043
`define RAMB36E2__INIT_29_SZ 256

`define RAMB36E2__INIT_2A    32'h00000044
`define RAMB36E2__INIT_2A_SZ 256

`define RAMB36E2__INIT_2B    32'h00000045
`define RAMB36E2__INIT_2B_SZ 256

`define RAMB36E2__INIT_2C    32'h00000046
`define RAMB36E2__INIT_2C_SZ 256

`define RAMB36E2__INIT_2D    32'h00000047
`define RAMB36E2__INIT_2D_SZ 256

`define RAMB36E2__INIT_2E    32'h00000048
`define RAMB36E2__INIT_2E_SZ 256

`define RAMB36E2__INIT_2F    32'h00000049
`define RAMB36E2__INIT_2F_SZ 256

`define RAMB36E2__INIT_30    32'h0000004a
`define RAMB36E2__INIT_30_SZ 256

`define RAMB36E2__INIT_31    32'h0000004b
`define RAMB36E2__INIT_31_SZ 256

`define RAMB36E2__INIT_32    32'h0000004c
`define RAMB36E2__INIT_32_SZ 256

`define RAMB36E2__INIT_33    32'h0000004d
`define RAMB36E2__INIT_33_SZ 256

`define RAMB36E2__INIT_34    32'h0000004e
`define RAMB36E2__INIT_34_SZ 256

`define RAMB36E2__INIT_35    32'h0000004f
`define RAMB36E2__INIT_35_SZ 256

`define RAMB36E2__INIT_36    32'h00000050
`define RAMB36E2__INIT_36_SZ 256

`define RAMB36E2__INIT_37    32'h00000051
`define RAMB36E2__INIT_37_SZ 256

`define RAMB36E2__INIT_38    32'h00000052
`define RAMB36E2__INIT_38_SZ 256

`define RAMB36E2__INIT_39    32'h00000053
`define RAMB36E2__INIT_39_SZ 256

`define RAMB36E2__INIT_3A    32'h00000054
`define RAMB36E2__INIT_3A_SZ 256

`define RAMB36E2__INIT_3B    32'h00000055
`define RAMB36E2__INIT_3B_SZ 256

`define RAMB36E2__INIT_3C    32'h00000056
`define RAMB36E2__INIT_3C_SZ 256

`define RAMB36E2__INIT_3D    32'h00000057
`define RAMB36E2__INIT_3D_SZ 256

`define RAMB36E2__INIT_3E    32'h00000058
`define RAMB36E2__INIT_3E_SZ 256

`define RAMB36E2__INIT_3F    32'h00000059
`define RAMB36E2__INIT_3F_SZ 256

`define RAMB36E2__INIT_40    32'h0000005a
`define RAMB36E2__INIT_40_SZ 256

`define RAMB36E2__INIT_41    32'h0000005b
`define RAMB36E2__INIT_41_SZ 256

`define RAMB36E2__INIT_42    32'h0000005c
`define RAMB36E2__INIT_42_SZ 256

`define RAMB36E2__INIT_43    32'h0000005d
`define RAMB36E2__INIT_43_SZ 256

`define RAMB36E2__INIT_44    32'h0000005e
`define RAMB36E2__INIT_44_SZ 256

`define RAMB36E2__INIT_45    32'h0000005f
`define RAMB36E2__INIT_45_SZ 256

`define RAMB36E2__INIT_46    32'h00000060
`define RAMB36E2__INIT_46_SZ 256

`define RAMB36E2__INIT_47    32'h00000061
`define RAMB36E2__INIT_47_SZ 256

`define RAMB36E2__INIT_48    32'h00000062
`define RAMB36E2__INIT_48_SZ 256

`define RAMB36E2__INIT_49    32'h00000063
`define RAMB36E2__INIT_49_SZ 256

`define RAMB36E2__INIT_4A    32'h00000064
`define RAMB36E2__INIT_4A_SZ 256

`define RAMB36E2__INIT_4B    32'h00000065
`define RAMB36E2__INIT_4B_SZ 256

`define RAMB36E2__INIT_4C    32'h00000066
`define RAMB36E2__INIT_4C_SZ 256

`define RAMB36E2__INIT_4D    32'h00000067
`define RAMB36E2__INIT_4D_SZ 256

`define RAMB36E2__INIT_4E    32'h00000068
`define RAMB36E2__INIT_4E_SZ 256

`define RAMB36E2__INIT_4F    32'h00000069
`define RAMB36E2__INIT_4F_SZ 256

`define RAMB36E2__INIT_50    32'h0000006a
`define RAMB36E2__INIT_50_SZ 256

`define RAMB36E2__INIT_51    32'h0000006b
`define RAMB36E2__INIT_51_SZ 256

`define RAMB36E2__INIT_52    32'h0000006c
`define RAMB36E2__INIT_52_SZ 256

`define RAMB36E2__INIT_53    32'h0000006d
`define RAMB36E2__INIT_53_SZ 256

`define RAMB36E2__INIT_54    32'h0000006e
`define RAMB36E2__INIT_54_SZ 256

`define RAMB36E2__INIT_55    32'h0000006f
`define RAMB36E2__INIT_55_SZ 256

`define RAMB36E2__INIT_56    32'h00000070
`define RAMB36E2__INIT_56_SZ 256

`define RAMB36E2__INIT_57    32'h00000071
`define RAMB36E2__INIT_57_SZ 256

`define RAMB36E2__INIT_58    32'h00000072
`define RAMB36E2__INIT_58_SZ 256

`define RAMB36E2__INIT_59    32'h00000073
`define RAMB36E2__INIT_59_SZ 256

`define RAMB36E2__INIT_5A    32'h00000074
`define RAMB36E2__INIT_5A_SZ 256

`define RAMB36E2__INIT_5B    32'h00000075
`define RAMB36E2__INIT_5B_SZ 256

`define RAMB36E2__INIT_5C    32'h00000076
`define RAMB36E2__INIT_5C_SZ 256

`define RAMB36E2__INIT_5D    32'h00000077
`define RAMB36E2__INIT_5D_SZ 256

`define RAMB36E2__INIT_5E    32'h00000078
`define RAMB36E2__INIT_5E_SZ 256

`define RAMB36E2__INIT_5F    32'h00000079
`define RAMB36E2__INIT_5F_SZ 256

`define RAMB36E2__INIT_60    32'h0000007a
`define RAMB36E2__INIT_60_SZ 256

`define RAMB36E2__INIT_61    32'h0000007b
`define RAMB36E2__INIT_61_SZ 256

`define RAMB36E2__INIT_62    32'h0000007c
`define RAMB36E2__INIT_62_SZ 256

`define RAMB36E2__INIT_63    32'h0000007d
`define RAMB36E2__INIT_63_SZ 256

`define RAMB36E2__INIT_64    32'h0000007e
`define RAMB36E2__INIT_64_SZ 256

`define RAMB36E2__INIT_65    32'h0000007f
`define RAMB36E2__INIT_65_SZ 256

`define RAMB36E2__INIT_66    32'h00000080
`define RAMB36E2__INIT_66_SZ 256

`define RAMB36E2__INIT_67    32'h00000081
`define RAMB36E2__INIT_67_SZ 256

`define RAMB36E2__INIT_68    32'h00000082
`define RAMB36E2__INIT_68_SZ 256

`define RAMB36E2__INIT_69    32'h00000083
`define RAMB36E2__INIT_69_SZ 256

`define RAMB36E2__INIT_6A    32'h00000084
`define RAMB36E2__INIT_6A_SZ 256

`define RAMB36E2__INIT_6B    32'h00000085
`define RAMB36E2__INIT_6B_SZ 256

`define RAMB36E2__INIT_6C    32'h00000086
`define RAMB36E2__INIT_6C_SZ 256

`define RAMB36E2__INIT_6D    32'h00000087
`define RAMB36E2__INIT_6D_SZ 256

`define RAMB36E2__INIT_6E    32'h00000088
`define RAMB36E2__INIT_6E_SZ 256

`define RAMB36E2__INIT_6F    32'h00000089
`define RAMB36E2__INIT_6F_SZ 256

`define RAMB36E2__INIT_70    32'h0000008a
`define RAMB36E2__INIT_70_SZ 256

`define RAMB36E2__INIT_71    32'h0000008b
`define RAMB36E2__INIT_71_SZ 256

`define RAMB36E2__INIT_72    32'h0000008c
`define RAMB36E2__INIT_72_SZ 256

`define RAMB36E2__INIT_73    32'h0000008d
`define RAMB36E2__INIT_73_SZ 256

`define RAMB36E2__INIT_74    32'h0000008e
`define RAMB36E2__INIT_74_SZ 256

`define RAMB36E2__INIT_75    32'h0000008f
`define RAMB36E2__INIT_75_SZ 256

`define RAMB36E2__INIT_76    32'h00000090
`define RAMB36E2__INIT_76_SZ 256

`define RAMB36E2__INIT_77    32'h00000091
`define RAMB36E2__INIT_77_SZ 256

`define RAMB36E2__INIT_78    32'h00000092
`define RAMB36E2__INIT_78_SZ 256

`define RAMB36E2__INIT_79    32'h00000093
`define RAMB36E2__INIT_79_SZ 256

`define RAMB36E2__INIT_7A    32'h00000094
`define RAMB36E2__INIT_7A_SZ 256

`define RAMB36E2__INIT_7B    32'h00000095
`define RAMB36E2__INIT_7B_SZ 256

`define RAMB36E2__INIT_7C    32'h00000096
`define RAMB36E2__INIT_7C_SZ 256

`define RAMB36E2__INIT_7D    32'h00000097
`define RAMB36E2__INIT_7D_SZ 256

`define RAMB36E2__INIT_7E    32'h00000098
`define RAMB36E2__INIT_7E_SZ 256

`define RAMB36E2__INIT_7F    32'h00000099
`define RAMB36E2__INIT_7F_SZ 256

`define RAMB36E2__INIT_A    32'h0000009a
`define RAMB36E2__INIT_A_SZ 36

`define RAMB36E2__INIT_B    32'h0000009b
`define RAMB36E2__INIT_B_SZ 36

`define RAMB36E2__INIT_FILE    32'h0000009c
`define RAMB36E2__INIT_FILE_SZ 32

`define RAMB36E2__IS_CLKARDCLK_INVERTED    32'h0000009d
`define RAMB36E2__IS_CLKARDCLK_INVERTED_SZ 1

`define RAMB36E2__IS_CLKBWRCLK_INVERTED    32'h0000009e
`define RAMB36E2__IS_CLKBWRCLK_INVERTED_SZ 1

`define RAMB36E2__IS_ENARDEN_INVERTED    32'h0000009f
`define RAMB36E2__IS_ENARDEN_INVERTED_SZ 1

`define RAMB36E2__IS_ENBWREN_INVERTED    32'h000000a0
`define RAMB36E2__IS_ENBWREN_INVERTED_SZ 1

`define RAMB36E2__IS_RSTRAMARSTRAM_INVERTED    32'h000000a1
`define RAMB36E2__IS_RSTRAMARSTRAM_INVERTED_SZ 1

`define RAMB36E2__IS_RSTRAMB_INVERTED    32'h000000a2
`define RAMB36E2__IS_RSTRAMB_INVERTED_SZ 1

`define RAMB36E2__IS_RSTREGARSTREG_INVERTED    32'h000000a3
`define RAMB36E2__IS_RSTREGARSTREG_INVERTED_SZ 1

`define RAMB36E2__IS_RSTREGB_INVERTED    32'h000000a4
`define RAMB36E2__IS_RSTREGB_INVERTED_SZ 1

`define RAMB36E2__RDADDRCHANGEA    32'h000000a5
`define RAMB36E2__RDADDRCHANGEA_SZ 40

`define RAMB36E2__RDADDRCHANGEB    32'h000000a6
`define RAMB36E2__RDADDRCHANGEB_SZ 40

`define RAMB36E2__READ_WIDTH_A    32'h000000a7
`define RAMB36E2__READ_WIDTH_A_SZ 32

`define RAMB36E2__READ_WIDTH_B    32'h000000a8
`define RAMB36E2__READ_WIDTH_B_SZ 32

`define RAMB36E2__RSTREG_PRIORITY_A    32'h000000a9
`define RAMB36E2__RSTREG_PRIORITY_A_SZ 48

`define RAMB36E2__RSTREG_PRIORITY_B    32'h000000aa
`define RAMB36E2__RSTREG_PRIORITY_B_SZ 48

`define RAMB36E2__SIM_COLLISION_CHECK    32'h000000ab
`define RAMB36E2__SIM_COLLISION_CHECK_SZ 120

`define RAMB36E2__SLEEP_ASYNC    32'h000000ac
`define RAMB36E2__SLEEP_ASYNC_SZ 40

`define RAMB36E2__SRVAL_A    32'h000000ad
`define RAMB36E2__SRVAL_A_SZ 36

`define RAMB36E2__SRVAL_B    32'h000000ae
`define RAMB36E2__SRVAL_B_SZ 36

`define RAMB36E2__WRITE_MODE_A    32'h000000af
`define RAMB36E2__WRITE_MODE_A_SZ 88

`define RAMB36E2__WRITE_MODE_B    32'h000000b0
`define RAMB36E2__WRITE_MODE_B_SZ 88

`define RAMB36E2__WRITE_WIDTH_A    32'h000000b1
`define RAMB36E2__WRITE_WIDTH_A_SZ 32

`define RAMB36E2__WRITE_WIDTH_B    32'h000000b2
`define RAMB36E2__WRITE_WIDTH_B_SZ 32

`endif  // B_RAMB36E2_DEFINES_VH