`include "B_VDU_defines.vh"

reg [`VDU_DATA_SZ-1:0] ATTR [0:`VDU_ADDR_N-1];
reg [`VDU__CORE_CODING_STANDARD_SZ:1] CORE_CODING_STANDARD_REG = CORE_CODING_STANDARD;
reg [`VDU__CORE_COLOR_DEPTH_SZ-1:0] CORE_COLOR_DEPTH_REG = CORE_COLOR_DEPTH;
reg [`VDU__CORE_COLOR_FORMAT_SZ-1:0] CORE_COLOR_FORMAT_REG = CORE_COLOR_FORMAT;
reg [`VDU__CORE_FRAME_PER_SECOND_SZ-1:0] CORE_FRAME_PER_SECOND_REG = CORE_FRAME_PER_SECOND;
reg [`VDU__CORE_FRAME_TYPE_SZ:1] CORE_FRAME_TYPE_REG = CORE_FRAME_TYPE;
real CORE_FREQUENCY_REG = CORE_FREQUENCY;
reg [`VDU__CORE_NO_OF_STREAMS_SZ-1:0] CORE_NO_OF_STREAMS_REG = CORE_NO_OF_STREAMS;
reg [`VDU__CORE_RESOLUTION_SZ:1] CORE_RESOLUTION_REG = CORE_RESOLUTION;

initial begin
  ATTR[`VDU__CORE_CODING_STANDARD] = CORE_CODING_STANDARD;
  ATTR[`VDU__CORE_COLOR_DEPTH] = CORE_COLOR_DEPTH;
  ATTR[`VDU__CORE_COLOR_FORMAT] = CORE_COLOR_FORMAT;
  ATTR[`VDU__CORE_FRAME_PER_SECOND] = CORE_FRAME_PER_SECOND;
  ATTR[`VDU__CORE_FRAME_TYPE] = CORE_FRAME_TYPE;
  ATTR[`VDU__CORE_FREQUENCY] = $realtobits(CORE_FREQUENCY);
  ATTR[`VDU__CORE_NO_OF_STREAMS] = CORE_NO_OF_STREAMS;
  ATTR[`VDU__CORE_RESOLUTION] = CORE_RESOLUTION;
end

always @(trig_attr) begin
  CORE_CODING_STANDARD_REG = ATTR[`VDU__CORE_CODING_STANDARD];
  CORE_COLOR_DEPTH_REG = ATTR[`VDU__CORE_COLOR_DEPTH];
  CORE_COLOR_FORMAT_REG = ATTR[`VDU__CORE_COLOR_FORMAT];
  CORE_FRAME_PER_SECOND_REG = ATTR[`VDU__CORE_FRAME_PER_SECOND];
  CORE_FRAME_TYPE_REG = ATTR[`VDU__CORE_FRAME_TYPE];
  CORE_FREQUENCY_REG = $bitstoreal(ATTR[`VDU__CORE_FREQUENCY]);
  CORE_NO_OF_STREAMS_REG = ATTR[`VDU__CORE_NO_OF_STREAMS];
  CORE_RESOLUTION_REG = ATTR[`VDU__CORE_RESOLUTION];
end

// procedures to override, read attribute values

task write_attr;
  input  [`VDU_ADDR_SZ-1:0] addr;
  input  [`VDU_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`VDU_DATA_SZ-1:0] read_attr;
  input  [`VDU_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
