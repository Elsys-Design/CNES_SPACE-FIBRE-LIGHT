library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.data_link_lib.all;

entity data_link is
  generic(
    G_VC_NUM           : integer := 8                                                  --! Number of virtual channel
    );
  port(
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- Network layer AXI-Stream TX interface
    AXIS_ACLK_TX_DL        : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_TX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_TX_DL       : in  vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_TX_DL       : in  vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_TX_DL       : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_TX_DL      : in  std_logic_vector(G_VC_NUM downto 0);
    -- Network layer RX interface
    AXIS_ACLK_RX_DL        : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_RX_DL      : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_RX_DL       : out vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_RX_DL       : out vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_RX_DL       : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_RX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    -- Lane layer TX interface
    DATA_TX_PPL            : out  std_logic_vector(31 downto 00);     --! Data parallel to be send from Data-Link Layer
    CAPABILITY_TX_PPL      : out  std_logic_vector(07 downto 00);     --! Capability send on TX link in INIT3 control word
    NEW_DATA_TX_PPL        : out  std_logic;                          --! Flag to write data in FIFO TX
    VALID_K_CHARAC_TX_PPL  : out  std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TX_PPL vector
    FIFO_TX_FULL_PPL       : in   std_logic;                          --! Flag full of the FIFO TX
    -- Lane layer RX interface
    FIFO_RX_RD_EN_PPL      : out  std_logic;                          --! Flag to read data in FIFO RX
    DATA_RX_PPL            : in   std_logic_vector(31 downto 00);     --! Data parallel to be received to Data-Link Layer
    FIFO_RX_EMPTY_PPL      : in   std_logic;                          --! Flag EMPTY of the FIFO RX
    FIFO_RX_DATA_VALID_PPL : in   std_logic;                          --! Flag DATA_VALID of the FIFO RX
    VALID_K_CHARAC_RX_PPL  : in   std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TR_PPL vector
    FAR_END_CAPA_DL        : in   std_logic_vector(07 downto 00);     --! Capability field receive in INIT3 control word
    -- MIB  parameters interface
    INTERFACE_RESET_DL     : in std_logic;                            --! Reset the link and all configuration register of the Data Link layer
    LINK_RESET_DL          : in std_logic;                            --! Reset the link
    NACK_RST_EN_DL         : in std_logic;                            --! Enable automatic link reset on NACK reception
    NACK_RST_MODE_DL       : in std_logic;                            --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
    PAUSE_VC_DL            : in std_logic_vector(G_VC_NUM downto 0);         --! Pause the corresponding virtual channel after the end of current transmission
    CONTINUOUS_VC_DL       : in std_logic_vector(G_VC_NUM-1 downto 0);         --! Enable the corresponding virtual channel continuous mode   
    -- MIB  status interface
    SEQ_NUMBER_TX_DL        : out std_logic_vector(G_VC_NUM-1 downto 0);       --! SEQ_NUMBER in transmission
    SEQ_NUMBER_RX_DL        : out std_logic_vector(G_VC_NUM-1 downto 0);       --! SEQ_NUMBER in reception
    CREDIT_VC_DL            : out std_logic_vector(G_VC_NUM-1 downto 0);       --! Indicates if each corresponding far-end input buffer has credit
    FCT_CREDIT_OVERFLOW_DL  : out std_logic_vector(G_VC_NUM-1 downto 0);       --! Indicates overflow of each corresponding input buffer
    CRC_LONG_ERROR_DL       : out std_logic;                          --! CRC long error
    CRC_SHORT_ERROR_DL      : out std_logic;                          --! CRC short error
    FRAME_ERROR_DL          : out std_logic;                          --! Frame error
    SEQUENCE_ERROR_DL       : out std_logic;                          --! Sequence error
    FAR_END_LINK_RESET_DL   : out std_logic;                          --! Far-end link reset status
    FRAME_FINISHED_DL       : out std_logic_vector(G_VC_NUM downto 0);       --! Indicates that corresponding channel finished emitting a frame
    FRAME_TX_DL             : out std_logic_vector(G_VC_NUM downto 0);       --! Indicates that corresponding channel is emitting a frame
    DATA_COUNTER_TX_DL      : out std_logic_vector(6 downto 0);       --! Indicate the number of data transmitted in last frame emitted
    DATA_COUNTER_RX_DL      : out std_logic_vector(6 downto 0);       --! Indicate the number of data received in last frame received
    ACK_COUNTER_TX_DL       : out  std_logic_vector(2 downto 0);      --! ACK counter TX
    NACK_COUNTER_TX_DL      : out  std_logic_vector(2 downto 0);      --! NACK counter TX
    FCT_COUNTER_TX_DL       : out  std_logic_vector(3 downto 0);      --! FCT counter TX
    ACK_COUNTER_RX_DL       : out  std_logic_vector(2 downto 0);      --! ACK counter RX
    NACK_COUNTER_RX_DL      : out  std_logic_vector(2 downto 0);      --! NACK counter RX
    FCT_COUNTER_RX_DL       : out  std_logic_vector(3 downto 0);      --! FCT counter RX
    FULL_COUNTER_RX_DL      : out  std_logic_vector(1 downto 0);      --! FULL counter RX
    RETRY_COUNTER_RX_DL     : out  std_logic_vector(1 downto 0);      --! RETRY counter RX
    CURRENT_TIME_SLOT_DL    : out  std_logic_vector(7 downto 0)       --! Current time slot
  );
end data_link;

architecture Behavioral of data_link is
  -- Déclaration des composants
  component data_out_buff is
    port (
      RST_N                 : in  std_logic;
      CLK                   : in  std_logic;
      LINK_RESET            : in std_logic;
      S_AXIS_ACLK           : in std_logic;
      S_AXIS_TREADY         : out std_logic;
      S_AXIS_TDATA          : in std_logic_vector(C_DATA_LENGTH-1 downto 0);
      S_AXIS_TUSER          : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      S_AXIS_TLAST          : in std_logic;
      S_AXIS_TVALID         : in std_logic;
      VC_READY_DOBUF        : out  std_logic;
      DATA_DOBUF            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DOBUF  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      DATA_VALID_DOBUF      : out  std_logic;
      END_PACKET_DOBUF      : out  std_logic;
      VC_RD_EN_DMAC         : in   std_logic;
      M_VAL_DDES            : in std_logic_vector(C_M_SIZE-1 downto 0);
      FCT_FAR_END_DDES      : in std_logic;
      LANE_ACTIVE_ST_PPL    : in std_logic;
      FCT_CC_OVF_DOBUF      : out std_logic;
      VC_CONT_MODE_MIB      : in std_logic
    );
  end component;

  component data_mac is
    generic(
      G_VC_NUM           : integer := 8
    );
    port (
      RST_N              : in  std_logic;
      CLK                : in  std_logic;
      REQ_ACK_DERRM       : in  std_logic;
      REQ_NACK_DERRM      : in  std_logic;
      TRANS_POL_FLG_DERRM : in  std_logic;
      REQ_ACK_DONE_DMAC   : out std_logic;
      REQ_FCT_DIBUF       : in  std_logic_vector(G_VC_NUM-1 downto 0);
      REQ_FCT_DONE_DIBUF  : out std_logic_vector(G_VC_NUM-1 downto 0);
      VC_READY_DOBUF      : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_DATA_DOBUF       : in  vc_data_array(G_VC_NUM-1 downto 0);
      VC_DATA_VALID_DOBUF : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_RD_EN_DMAC       : out  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_PAUSE_MIB        : in  std_logic_vector(G_VC_NUM-1 downto 0);
      VC_END_EMISSION_MIB : out std_logic_vector(G_VC_NUM-1 downto 0);
      VC_RUN_EMISSION_MIB : out std_logic_vector(G_VC_NUM-1 downto 0);
      DATA_DMAC            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);
      NEW_WORD_DMAC        : out std_logic;
      NEW_PACKET_DMAC      : out std_logic;
      END_PACKET_DMAC      : out std_logic;
      TYPE_FRAME_DMAC      : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      VIRTUAL_CHANNEL_DMAC : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_TYPE_DMAC         : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_CHANNEL_DMAC      : out std_logic_vector(G_VC_NUM-1 downto 0);
      BC_STATUS_DMAC       : out std_logic_vector(2-1 downto 0);
      MULT_CHANNEL_DMAC    : out std_logic_vector(G_VC_NUM-1 downto 0);
      TRANS_POL_FLG_DMAC   : out std_logic;
      READY_DENC           : in std_logic
    );
  end component;

  component data_encpasulation is
    generic (
        G_VC_NUM : integer := 8
    );
    port (
      RST_N                 : in  std_logic;
      CLK                   : in  std_logic;
      DATA_DMAC             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      NEW_WORD_DMAC         : in  std_logic;
      NEW_PACKET_DMAC       : in  std_logic;
      END_PACKET_DMAC       : in  std_logic;
      TYPE_FRAME_DMAC       : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      VIRTUAL_CHANNEL_DMAC  : in std_logic_vector (G_VC_NUM-1 downto 0);
      BC_TYPE_DMAC          : in std_logic_vector (G_VC_NUM-1 downto 0);
      BC_CHANNEL_DMAC       : in std_logic_vector (G_VC_NUM-1 downto 0);
      BC_STATUS_DMAC        : in std_logic_vector (2-1 downto 0);
      MULT_CHANNEL_DMAC     : in std_logic_vector (G_VC_NUM-1 downto 0);
      READY_DENC            : out std_logic;
      NEW_WORD_DENC         : out  std_logic;
      DATA_DENC             : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DENC   : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      TYPE_FRAME_DENC       : out  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      END_FRAME_DENC        : out  std_logic
    );
  end component;

  component data_seq_compute is
    port (
      RST_N                 : in  std_logic;
      CLK                   : in  std_logic;
      NEW_WORD_DENC         : in  std_logic;
      DATA_DENC             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DENC   : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      TYPE_FRAME_DENC       : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      END_FRAME_DENC        : in  std_logic;
      NEW_WORD_DSCOM        : out  std_logic;
      DATA_DSCOM            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DSCOM  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      TYPE_FRAME_DSCOM      : out  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      END_FRAME_DSCOM       : out  std_logic
    );
  end component;

  component data_crc_compute is
    port (
      RST_N                 : in  std_logic;
      CLK                   : in  std_logic;
      NEW_WORD_DSCOM        : in  std_logic;
      DATA_DSCOM            : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      VALID_K_CHARAC_DSCOM  : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      TYPE_FRAME_DSCOM      : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
      END_FRAME_DSCOM       : in  std_logic;
      FIFO_FULL_TX_LANE     : in  std_logic;
      VALID_K_CHARAC_DCCOM  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
      DATA_DCCOM            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);
      NEW_WORD_DCCOM        : out  std_logic
    );
  end component;

  -- Signaux internes
  signal link_reset            : std_logic;
  signal lane_active_st_ppl    : std_logic;
  -- MIB 
  signal vc_cont_mode_mib      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal vc_end_emission_mib  : std_logic_vector(G_VC_NUM-1 downto 0);
  signal vc_run_emission_mib  : std_logic_vector(G_VC_NUM-1 downto 0);
  signal vc_pause_mib         : std_logic_vector(G_VC_NUM-1 downto 0);
  -- Input Buffer
  signal req_fct_dibuf        : std_logic_vector(G_VC_NUM-1 downto 0);
  signal req_fct_done_dibuf   : std_logic_vector(G_VC_NUM-1 downto 0);
  -- Desencapsulation
  signal m_val_ddes            : vc_mult_array(G_VC_NUM-1 downto 0);
  signal fct_far_end_ddes      : std_logic_vector(G_VC_NUM-1 downto 0);
  -- Error Management
  signal req_ack_derrm        : std_logic;
  signal req_nack_derrm       : std_logic;
  signal trans_pol_flg_derrm  : std_logic;
  -- Output Buffer 
  signal vc_ready_dobuf        : std_logic_vector(G_VC_NUM-1 downto 0);
  signal vc_data_dobuf            : vc_data_array(G_VC_NUM-1 downto 0);
  signal valid_k_charac_dobuf  : vc_k_array(G_VC_NUM-1 downto 0);
  signal vc_data_valid_dobuf      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal end_packet_dobuf      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal fct_cc_ovf_dobuf      : std_logic_vector(G_VC_NUM-1 downto 0);
  -- Medium Acces Controller
  signal data_dmac             : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal new_word_dmac         : std_logic;
  signal new_packet_dmac      : std_logic;
  signal end_packet_dmac      : std_logic;
  signal type_frame_dmac      : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal virtual_channel_dmaC : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_type_dmac         : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_channel_dmac      : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_status_dmac       : std_logic_vector(2-1 downto 0);
  signal mult_channel_dmac    : std_logic_vector(G_VC_NUM-1 downto 0);
  signal trans_pol_flg_dmac   : std_logic;
  signal req_ack_done_dmac    : std_logic;
  signal vc_rd_en_dmac        : std_logic_vector(G_VC_NUM-1 downto 0);
  -- Encapsulation
  signal new_word_denc        : std_logic;
  signal data_denc            : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_denc  : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal type_frame_denc      : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal end_frame_denc       : std_logic;
  signal ready_denc           : std_logic;
  -- SEQ compute
  signal new_word_dscom       : std_logic;
  signal data_dscom           : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dscom : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal type_frame_dscom     : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal end_frame_dscom      : std_logic;
  -- CRC comppute 
  signal valid_k_charac_dccom : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal data_dccom           : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal new_word_dccom       : std_logic;

begin
  
  gen_data_out_buff: for i in 0 to G_VC_NUM-1 generate
    inst_data_out_buff: data_out_buff
      port map (
        RST_N                 => rst_n,
        CLK                   => clk,
        LINK_RESET            => link_reset,
        S_AXIS_ACLK           => axis_aclk_tx_dl(i),
        S_AXIS_TREADY         => axis_tready_tx_dl(i),
        S_AXIS_TDATA          => axis_tdata_tx_dl(i),
        S_AXIS_TUSER          => axis_tuser_tx_dl(i),
        S_AXIS_TLAST          => axis_tlast_tx_dl(i),
        S_AXIS_TVALID         => axis_tvalid_tx_dl(i),
        VC_READY_DOBUF        => vc_ready_dobuf(i),
        DATA_DOBUF            => vc_data_dobuf(i),
        VALID_K_CHARAC_DOBUF  => valid_k_charac_dobuf(i),
        DATA_VALID_DOBUF      => vc_data_valid_dobuf(i),
        END_PACKET_DOBUF      => end_packet_dobuf(i),
        VC_RD_EN_DMAC         => vc_rd_en_dmac(i),
        M_VAL_DDES            => m_val_ddes(i),
        FCT_FAR_END_DDES      => fct_far_end_ddes(i),
        LANE_ACTIVE_ST_PPL    => lane_active_st_ppl,
        FCT_CC_OVF_DOBUF      => fct_cc_ovf_dobuf(i),
        VC_CONT_MODE_MIB      => vc_cont_mode_mib(i)
      );
  end generate;

  inst_data_mac: data_mac
    generic map (
      G_VC_NUM => g_vc_num
    )
    port map (
      RST_N                => rst_n,
      CLK                  => clk,
      REQ_ACK_DERRM        => req_ack_derrm,
      REQ_NACK_DERRM       => req_nack_derrm,
      TRANS_POL_FLG_DERRM  => trans_pol_flg_derrm,
      REQ_ACK_DONE_DMAC    => req_ack_done_dmac,
      REQ_FCT_DONE_DIBUF   => req_fct_done_dibuf,
      REQ_FCT_DIBUF        => req_fct_dibuf,
      VC_READY_DOBUF       => vc_ready_dobuf,
      VC_DATA_DOBUF        => vc_data_dobuf,
      VC_DATA_VALID_DOBUF  => vc_data_valid_dobuf,
      VC_RD_EN_DMAC        => vc_rd_en_dmac,
      VC_PAUSE_MIB         => vc_pause_mib,
      VC_END_EMISSION_MIB  => vc_end_emission_mib,
      VC_RUN_EMISSION_MIB  => vc_run_emission_mib,
      DATA_DMAC            => data_dmac,
      NEW_WORD_DMAC        => new_word_dmac,
      NEW_PACKET_DMAC      => new_packet_dmac,
      END_PACKET_DMAC      => end_packet_dmac,
      TYPE_FRAME_DMAC      => type_frame_dmac,
      VIRTUAL_CHANNEL_DMAC => virtual_channel_dmac,
      BC_TYPE_DMAC         => bc_type_dmac,
      BC_CHANNEL_DMAC      => bc_channel_dmac,
      BC_STATUS_DMAC       => bc_status_dmac,
      MULT_CHANNEL_DMAC    => mult_channel_dmac,
      TRANS_POL_FLG_DMAC   => trans_pol_flg_dmac,
      READY_DENC           => ready_denc
    );

  inst_data_encpasulation: data_encpasulation
    generic map (
      G_VC_NUM => g_vc_num
    )
    port map (
      RST_N                 => rst_n,
      CLK                   => clk,
      DATA_DMAC             => data_dmac,
      NEW_WORD_DMAC         => new_word_dmac,
      NEW_PACKET_DMAC       => new_packet_dmac,
      END_PACKET_DMAC       => end_packet_dmac,
      TYPE_FRAME_DMAC       => type_frame_dmac,
      VIRTUAL_CHANNEL_DMAC  => virtual_channel_dmac,
      BC_TYPE_DMAC          => bc_type_dmac,
      BC_CHANNEL_DMAC       => bc_channel_dmac,
      BC_STATUS_DMAC        => bc_status_dmac,
      MULT_CHANNEL_DMAC     => mult_channel_dmac,
      READY_DENC            => ready_denc,
      NEW_WORD_DENC         => new_word_denc,
      DATA_DENC             => data_denc,
      VALID_K_CHARAC_DENC   => valid_k_charac_denc,
      TYPE_FRAME_DENC       => type_frame_denc,
      END_FRAME_DENC        => end_frame_denc
    );

  inst_data_seq_compute: data_seq_compute
    port map (
      RST_N                 => rst_n,
      CLK                   => clk,
      NEW_WORD_DENC         => new_word_denc,
      DATA_DENC             => data_denc,
      VALID_K_CHARAC_DENC   => valid_k_charac_denc,
      TYPE_FRAME_DENC       => type_frame_denc,
      END_FRAME_DENC        => end_frame_denc,
      NEW_WORD_DSCOM        => new_word_dscom,
      DATA_DSCOM            => data_dscom,
      VALID_K_CHARAC_DSCOM  => valid_k_charac_dscom,
      TYPE_FRAME_DSCOM      => type_frame_dscom,
      END_FRAME_DSCOM       => end_frame_dscom
    );

  inst_data_crc_compute: data_crc_compute
    port map (
      RST_N                 => rst_n,
      CLK                   => clk,
      NEW_WORD_DSCOM        => new_word_dscom,
      DATA_DSCOM            => data_dscom,
      VALID_K_CHARAC_DSCOM  => valid_k_charac_dscom,
      TYPE_FRAME_DSCOM      => type_frame_dscom,
      END_FRAME_DSCOM       => end_frame_dscom,
      FIFO_FULL_TX_LANE     => FIFO_TX_FULL_PPL,
      VALID_K_CHARAC_DCCOM  => valid_k_charac_dccom,
      DATA_DCCOM            => data_dccom,
      NEW_WORD_DCCOM        => new_word_dccom
    );

end Behavioral;
