// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC_NCRB_SSIT_DEFINES_VH
`else
`define B_NOC_NCRB_SSIT_DEFINES_VH

// Look-up table parameters
//

`define NOC_NCRB_SSIT_ADDR_N  9
`define NOC_NCRB_SSIT_ADDR_SZ 32
`define NOC_NCRB_SSIT_DATA_SZ 32

// Attribute addresses
//

`define NOC_NCRB_SSIT__REG_P0_0_VCA_TOKEN    32'h00000000
`define NOC_NCRB_SSIT__REG_P0_0_VCA_TOKEN_SZ 32

`define NOC_NCRB_SSIT__REG_P0_1_VCA_TOKEN    32'h00000001
`define NOC_NCRB_SSIT__REG_P0_1_VCA_TOKEN_SZ 32

`define NOC_NCRB_SSIT__REG_P0_R2W_EB_CTRL    32'h00000002
`define NOC_NCRB_SSIT__REG_P0_R2W_EB_CTRL_SZ 21

`define NOC_NCRB_SSIT__REG_P0_W2R_EB_CTRL    32'h00000003
`define NOC_NCRB_SSIT__REG_P0_W2R_EB_CTRL_SZ 21

`define NOC_NCRB_SSIT__REG_P1_0_VCA_TOKEN    32'h00000004
`define NOC_NCRB_SSIT__REG_P1_0_VCA_TOKEN_SZ 32

`define NOC_NCRB_SSIT__REG_P1_1_VCA_TOKEN    32'h00000005
`define NOC_NCRB_SSIT__REG_P1_1_VCA_TOKEN_SZ 32

`define NOC_NCRB_SSIT__REG_P1_R2W_EB_CTRL    32'h00000006
`define NOC_NCRB_SSIT__REG_P1_R2W_EB_CTRL_SZ 21

`define NOC_NCRB_SSIT__REG_P1_W2R_EB_CTRL    32'h00000007
`define NOC_NCRB_SSIT__REG_P1_W2R_EB_CTRL_SZ 21

`define NOC_NCRB_SSIT__REG_PIPE_MODE    32'h00000008
`define NOC_NCRB_SSIT__REG_PIPE_MODE_SZ 1

`endif  // B_NOC_NCRB_SSIT_DEFINES_VH