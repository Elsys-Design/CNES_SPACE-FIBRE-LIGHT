// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IDELAYE3_DEFINES_VH
`else
`define B_IDELAYE3_DEFINES_VH

// Look-up table parameters
//

`define IDELAYE3_ADDR_N  12
`define IDELAYE3_ADDR_SZ 32
`define IDELAYE3_DATA_SZ 152

// Attribute addresses
//

`define IDELAYE3__CASCADE    32'h00000000
`define IDELAYE3__CASCADE_SZ 96

`define IDELAYE3__DELAY_FORMAT    32'h00000001
`define IDELAYE3__DELAY_FORMAT_SZ 40

`define IDELAYE3__DELAY_SRC    32'h00000002
`define IDELAYE3__DELAY_SRC_SZ 56

`define IDELAYE3__DELAY_TYPE    32'h00000003
`define IDELAYE3__DELAY_TYPE_SZ 64

`define IDELAYE3__DELAY_VALUE    32'h00000004
`define IDELAYE3__DELAY_VALUE_SZ 32

`define IDELAYE3__IS_CLK_INVERTED    32'h00000005
`define IDELAYE3__IS_CLK_INVERTED_SZ 1

`define IDELAYE3__IS_RST_INVERTED    32'h00000006
`define IDELAYE3__IS_RST_INVERTED_SZ 1

`define IDELAYE3__LOOPBACK    32'h00000007
`define IDELAYE3__LOOPBACK_SZ 40

`define IDELAYE3__REFCLK_FREQUENCY    32'h00000008
`define IDELAYE3__REFCLK_FREQUENCY_SZ 64

`define IDELAYE3__SIM_DEVICE    32'h00000009
`define IDELAYE3__SIM_DEVICE_SZ 152

`define IDELAYE3__SIM_VERSION    32'h0000000a
`define IDELAYE3__SIM_VERSION_SZ 64

`define IDELAYE3__UPDATE_MODE    32'h0000000b
`define IDELAYE3__UPDATE_MODE_SZ 48

`endif  // B_IDELAYE3_DEFINES_VH