// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_X5PHIO_CMU_X32_DEFINES_VH
`else
`define B_X5PHIO_CMU_X32_DEFINES_VH

// Look-up table parameters
//

`define X5PHIO_CMU_X32_ADDR_N  61
`define X5PHIO_CMU_X32_ADDR_SZ 32
`define X5PHIO_CMU_X32_DATA_SZ 120

// Attribute addresses
//

`define X5PHIO_CMU_X32__ANATERM_NVAL    32'h00000000
`define X5PHIO_CMU_X32__ANATERM_NVAL_SZ 4

`define X5PHIO_CMU_X32__ANATERM_PVAL    32'h00000001
`define X5PHIO_CMU_X32__ANATERM_PVAL_SZ 4

`define X5PHIO_CMU_X32__ANATERM_SEL    32'h00000002
`define X5PHIO_CMU_X32__ANATERM_SEL_SZ 40

`define X5PHIO_CMU_X32__ATBMUX_SEL    32'h00000003
`define X5PHIO_CMU_X32__ATBMUX_SEL_SZ 12

`define X5PHIO_CMU_X32__ATB_PATH_SEL    32'h00000004
`define X5PHIO_CMU_X32__ATB_PATH_SEL_SZ 120

`define X5PHIO_CMU_X32__BYP_FREQ_DIV_S2P_CMU    32'h00000005
`define X5PHIO_CMU_X32__BYP_FREQ_DIV_S2P_CMU_SZ 40

`define X5PHIO_CMU_X32__BYP_FREQ_DIV_X5PLL    32'h00000006
`define X5PHIO_CMU_X32__BYP_FREQ_DIV_X5PLL_SZ 40

`define X5PHIO_CMU_X32__CALTX_RCAL_EN    32'h00000007
`define X5PHIO_CMU_X32__CALTX_RCAL_EN_SZ 40

`define X5PHIO_CMU_X32__CALTX_RCAL_VAL    32'h00000008
`define X5PHIO_CMU_X32__CALTX_RCAL_VAL_SZ 9

`define X5PHIO_CMU_X32__CMU_ADLY_BIAS    32'h00000009
`define X5PHIO_CMU_X32__CMU_ADLY_BIAS_SZ 3

`define X5PHIO_CMU_X32__CMU_APB_CLK_SEL    32'h0000000a
`define X5PHIO_CMU_X32__CMU_APB_CLK_SEL_SZ 104

`define X5PHIO_CMU_X32__CMU_CTLE_BIAS    32'h0000000b
`define X5PHIO_CMU_X32__CMU_CTLE_BIAS_SZ 5

`define X5PHIO_CMU_X32__CMU_D2C_BIAS    32'h0000000c
`define X5PHIO_CMU_X32__CMU_D2C_BIAS_SZ 3

`define X5PHIO_CMU_X32__CMU_DFE_BIAS    32'h0000000d
`define X5PHIO_CMU_X32__CMU_DFE_BIAS_SZ 11

`define X5PHIO_CMU_X32__CMU_LPRXBIAS_SEL    32'h0000000e
`define X5PHIO_CMU_X32__CMU_LPRXBIAS_SEL_SZ 5

`define X5PHIO_CMU_X32__CMU_NPI_CLK_SEL    32'h0000000f
`define X5PHIO_CMU_X32__CMU_NPI_CLK_SEL_SZ 104

`define X5PHIO_CMU_X32__CMU_RXBIAS_SPARE    32'h00000010
`define X5PHIO_CMU_X32__CMU_RXBIAS_SPARE_SZ 8

`define X5PHIO_CMU_X32__CMU_SRCH_ALGORITHM    32'h00000011
`define X5PHIO_CMU_X32__CMU_SRCH_ALGORITHM_SZ 48

`define X5PHIO_CMU_X32__CMU_TXBIAS_SEL    32'h00000012
`define X5PHIO_CMU_X32__CMU_TXBIAS_SEL_SZ 5

`define X5PHIO_CMU_X32__CMU_VREF_BIAS    32'h00000013
`define X5PHIO_CMU_X32__CMU_VREF_BIAS_SZ 7

`define X5PHIO_CMU_X32__DCI2LTCH_NCODE    32'h00000014
`define X5PHIO_CMU_X32__DCI2LTCH_NCODE_SZ 7

`define X5PHIO_CMU_X32__DCI2LTCH_PCODE    32'h00000015
`define X5PHIO_CMU_X32__DCI2LTCH_PCODE_SZ 7

`define X5PHIO_CMU_X32__DCIUPDATEMODE    32'h00000016
`define X5PHIO_CMU_X32__DCIUPDATEMODE_SZ 80

`define X5PHIO_CMU_X32__DCI_CASCADE_SEL    32'h00000017
`define X5PHIO_CMU_X32__DCI_CASCADE_SEL_SZ 2

`define X5PHIO_CMU_X32__DCI_CONFIG    32'h00000018
`define X5PHIO_CMU_X32__DCI_CONFIG_SZ 48

`define X5PHIO_CMU_X32__DCI_DEBUG_SEL    32'h00000019
`define X5PHIO_CMU_X32__DCI_DEBUG_SEL_SZ 16

`define X5PHIO_CMU_X32__DCI_FLTR_CTRL    32'h0000001a
`define X5PHIO_CMU_X32__DCI_FLTR_CTRL_SZ 4

`define X5PHIO_CMU_X32__DCI_ITER_SEL    32'h0000001b
`define X5PHIO_CMU_X32__DCI_ITER_SEL_SZ 88

`define X5PHIO_CMU_X32__DCI_LOCK_DIR    32'h0000001c
`define X5PHIO_CMU_X32__DCI_LOCK_DIR_SZ 40

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N0    32'h0000001d
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N0_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N1    32'h0000001e
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N1_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N2    32'h0000001f
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N2_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N3    32'h00000020
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N3_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N4    32'h00000021
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_N4_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P0    32'h00000022
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P0_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P1    32'h00000023
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P1_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P2    32'h00000024
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P2_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P3    32'h00000025
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P3_SZ 12

`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P4    32'h00000026
`define X5PHIO_CMU_X32__DCI_SCL_CTRL_P4_SZ 12

`define X5PHIO_CMU_X32__DCI_TYPE    32'h00000027
`define X5PHIO_CMU_X32__DCI_TYPE_SZ 6

`define X5PHIO_CMU_X32__DEBUG_CALTX_RCAL_EN    32'h00000028
`define X5PHIO_CMU_X32__DEBUG_CALTX_RCAL_EN_SZ 40

`define X5PHIO_CMU_X32__DEBUG_CALTX_RCAL_VAL    32'h00000029
`define X5PHIO_CMU_X32__DEBUG_CALTX_RCAL_VAL_SZ 9

`define X5PHIO_CMU_X32__DEBUG_DCI_LOCK_DIR    32'h0000002a
`define X5PHIO_CMU_X32__DEBUG_DCI_LOCK_DIR_SZ 40

`define X5PHIO_CMU_X32__DEBUG_RCAL_M_OVERRIDE    32'h0000002b
`define X5PHIO_CMU_X32__DEBUG_RCAL_M_OVERRIDE_SZ 40

`define X5PHIO_CMU_X32__DEBUG_VREF_APB_SEL    32'h0000002c
`define X5PHIO_CMU_X32__DEBUG_VREF_APB_SEL_SZ 40

`define X5PHIO_CMU_X32__DEBUG_VREF_MONITOR    32'h0000002d
`define X5PHIO_CMU_X32__DEBUG_VREF_MONITOR_SZ 40

`define X5PHIO_CMU_X32__EN_DCI    32'h0000002e
`define X5PHIO_CMU_X32__EN_DCI_SZ 40

`define X5PHIO_CMU_X32__EN_OUT_FLTR    32'h0000002f
`define X5PHIO_CMU_X32__EN_OUT_FLTR_SZ 40

`define X5PHIO_CMU_X32__RCAL_BUS    32'h00000030
`define X5PHIO_CMU_X32__RCAL_BUS_SZ 9

`define X5PHIO_CMU_X32__RCAL_ITER_SEL    32'h00000031
`define X5PHIO_CMU_X32__RCAL_ITER_SEL_SZ 96

`define X5PHIO_CMU_X32__RCAL_MODE    32'h00000032
`define X5PHIO_CMU_X32__RCAL_MODE_SZ 80

`define X5PHIO_CMU_X32__RCAL_M_OVERRIDE    32'h00000033
`define X5PHIO_CMU_X32__RCAL_M_OVERRIDE_SZ 40

`define X5PHIO_CMU_X32__RCAL_SCALE    32'h00000034
`define X5PHIO_CMU_X32__RCAL_SCALE_SZ 13

`define X5PHIO_CMU_X32__TST_EN    32'h00000035
`define X5PHIO_CMU_X32__TST_EN_SZ 40

`define X5PHIO_CMU_X32__VREF_0P3_CODE    32'h00000036
`define X5PHIO_CMU_X32__VREF_0P3_CODE_SZ 10

`define X5PHIO_CMU_X32__VREF_0P5_CODE    32'h00000037
`define X5PHIO_CMU_X32__VREF_0P5_CODE_SZ 10

`define X5PHIO_CMU_X32__VREF_0P75_CODE    32'h00000038
`define X5PHIO_CMU_X32__VREF_0P75_CODE_SZ 10

`define X5PHIO_CMU_X32__VREF_12P5_CODE    32'h00000039
`define X5PHIO_CMU_X32__VREF_12P5_CODE_SZ 10

`define X5PHIO_CMU_X32__VREF_16P7_CODE    32'h0000003a
`define X5PHIO_CMU_X32__VREF_16P7_CODE_SZ 10

`define X5PHIO_CMU_X32__VREF_MONITOR    32'h0000003b
`define X5PHIO_CMU_X32__VREF_MONITOR_SZ 40

`define X5PHIO_CMU_X32__WAIT_BYPASS    32'h0000003c
`define X5PHIO_CMU_X32__WAIT_BYPASS_SZ 40

`endif  // B_X5PHIO_CMU_X32_DEFINES_VH