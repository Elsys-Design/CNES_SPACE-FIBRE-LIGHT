// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTM_DUAL_DEFINES_VH
`else
`define B_GTM_DUAL_DEFINES_VH

// Look-up table parameters
//

`define GTM_DUAL_ADDR_N  363
`define GTM_DUAL_ADDR_SZ 32
`define GTM_DUAL_DATA_SZ 152

// Attribute addresses
//

`define GTM_DUAL__A_CFG    32'h00000000
`define GTM_DUAL__A_CFG_SZ 16

`define GTM_DUAL__A_SDM_DATA_CFG0    32'h00000001
`define GTM_DUAL__A_SDM_DATA_CFG0_SZ 16

`define GTM_DUAL__A_SDM_DATA_CFG1    32'h00000002
`define GTM_DUAL__A_SDM_DATA_CFG1_SZ 16

`define GTM_DUAL__BIAS_CFG0    32'h00000003
`define GTM_DUAL__BIAS_CFG0_SZ 16

`define GTM_DUAL__BIAS_CFG1    32'h00000004
`define GTM_DUAL__BIAS_CFG1_SZ 16

`define GTM_DUAL__BIAS_CFG2    32'h00000005
`define GTM_DUAL__BIAS_CFG2_SZ 16

`define GTM_DUAL__BIAS_CFG3    32'h00000006
`define GTM_DUAL__BIAS_CFG3_SZ 16

`define GTM_DUAL__BIAS_CFG4    32'h00000007
`define GTM_DUAL__BIAS_CFG4_SZ 16

`define GTM_DUAL__BIAS_CFG5    32'h00000008
`define GTM_DUAL__BIAS_CFG5_SZ 16

`define GTM_DUAL__BIAS_CFG6    32'h00000009
`define GTM_DUAL__BIAS_CFG6_SZ 16

`define GTM_DUAL__BIAS_CFG7    32'h0000000a
`define GTM_DUAL__BIAS_CFG7_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG0    32'h0000000b
`define GTM_DUAL__CH0_A_CH_CFG0_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG1    32'h0000000c
`define GTM_DUAL__CH0_A_CH_CFG1_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG2    32'h0000000d
`define GTM_DUAL__CH0_A_CH_CFG2_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG3    32'h0000000e
`define GTM_DUAL__CH0_A_CH_CFG3_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG4    32'h0000000f
`define GTM_DUAL__CH0_A_CH_CFG4_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG5    32'h00000010
`define GTM_DUAL__CH0_A_CH_CFG5_SZ 16

`define GTM_DUAL__CH0_A_CH_CFG6    32'h00000011
`define GTM_DUAL__CH0_A_CH_CFG6_SZ 16

`define GTM_DUAL__CH0_RST_LP_CFG0    32'h00000012
`define GTM_DUAL__CH0_RST_LP_CFG0_SZ 16

`define GTM_DUAL__CH0_RST_LP_CFG1    32'h00000013
`define GTM_DUAL__CH0_RST_LP_CFG1_SZ 16

`define GTM_DUAL__CH0_RST_LP_CFG2    32'h00000014
`define GTM_DUAL__CH0_RST_LP_CFG2_SZ 16

`define GTM_DUAL__CH0_RST_LP_CFG3    32'h00000015
`define GTM_DUAL__CH0_RST_LP_CFG3_SZ 16

`define GTM_DUAL__CH0_RST_LP_CFG4    32'h00000016
`define GTM_DUAL__CH0_RST_LP_CFG4_SZ 16

`define GTM_DUAL__CH0_RST_LP_ID_CFG0    32'h00000017
`define GTM_DUAL__CH0_RST_LP_ID_CFG0_SZ 16

`define GTM_DUAL__CH0_RST_LP_ID_CFG1    32'h00000018
`define GTM_DUAL__CH0_RST_LP_ID_CFG1_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG0    32'h00000019
`define GTM_DUAL__CH0_RST_TIME_CFG0_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG1    32'h0000001a
`define GTM_DUAL__CH0_RST_TIME_CFG1_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG2    32'h0000001b
`define GTM_DUAL__CH0_RST_TIME_CFG2_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG3    32'h0000001c
`define GTM_DUAL__CH0_RST_TIME_CFG3_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG4    32'h0000001d
`define GTM_DUAL__CH0_RST_TIME_CFG4_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG5    32'h0000001e
`define GTM_DUAL__CH0_RST_TIME_CFG5_SZ 16

`define GTM_DUAL__CH0_RST_TIME_CFG6    32'h0000001f
`define GTM_DUAL__CH0_RST_TIME_CFG6_SZ 16

`define GTM_DUAL__CH0_RX_ADC_CFG0    32'h00000020
`define GTM_DUAL__CH0_RX_ADC_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_ADC_CFG1    32'h00000021
`define GTM_DUAL__CH0_RX_ADC_CFG1_SZ 16

`define GTM_DUAL__CH0_RX_ANA_CFG0    32'h00000022
`define GTM_DUAL__CH0_RX_ANA_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_ANA_CFG1    32'h00000023
`define GTM_DUAL__CH0_RX_ANA_CFG1_SZ 16

`define GTM_DUAL__CH0_RX_ANA_CFG2    32'h00000024
`define GTM_DUAL__CH0_RX_ANA_CFG2_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG0A    32'h00000025
`define GTM_DUAL__CH0_RX_APT_CFG0A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG0B    32'h00000026
`define GTM_DUAL__CH0_RX_APT_CFG0B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG10A    32'h00000027
`define GTM_DUAL__CH0_RX_APT_CFG10A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG10B    32'h00000028
`define GTM_DUAL__CH0_RX_APT_CFG10B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG11A    32'h00000029
`define GTM_DUAL__CH0_RX_APT_CFG11A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG11B    32'h0000002a
`define GTM_DUAL__CH0_RX_APT_CFG11B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG12A    32'h0000002b
`define GTM_DUAL__CH0_RX_APT_CFG12A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG12B    32'h0000002c
`define GTM_DUAL__CH0_RX_APT_CFG12B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG13A    32'h0000002d
`define GTM_DUAL__CH0_RX_APT_CFG13A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG13B    32'h0000002e
`define GTM_DUAL__CH0_RX_APT_CFG13B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG14A    32'h0000002f
`define GTM_DUAL__CH0_RX_APT_CFG14A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG14B    32'h00000030
`define GTM_DUAL__CH0_RX_APT_CFG14B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG15A    32'h00000031
`define GTM_DUAL__CH0_RX_APT_CFG15A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG15B    32'h00000032
`define GTM_DUAL__CH0_RX_APT_CFG15B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG16A    32'h00000033
`define GTM_DUAL__CH0_RX_APT_CFG16A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG16B    32'h00000034
`define GTM_DUAL__CH0_RX_APT_CFG16B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG17A    32'h00000035
`define GTM_DUAL__CH0_RX_APT_CFG17A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG17B    32'h00000036
`define GTM_DUAL__CH0_RX_APT_CFG17B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG18A    32'h00000037
`define GTM_DUAL__CH0_RX_APT_CFG18A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG18B    32'h00000038
`define GTM_DUAL__CH0_RX_APT_CFG18B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG19A    32'h00000039
`define GTM_DUAL__CH0_RX_APT_CFG19A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG19B    32'h0000003a
`define GTM_DUAL__CH0_RX_APT_CFG19B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG1A    32'h0000003b
`define GTM_DUAL__CH0_RX_APT_CFG1A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG1B    32'h0000003c
`define GTM_DUAL__CH0_RX_APT_CFG1B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG20A    32'h0000003d
`define GTM_DUAL__CH0_RX_APT_CFG20A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG20B    32'h0000003e
`define GTM_DUAL__CH0_RX_APT_CFG20B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG21A    32'h0000003f
`define GTM_DUAL__CH0_RX_APT_CFG21A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG21B    32'h00000040
`define GTM_DUAL__CH0_RX_APT_CFG21B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG22A    32'h00000041
`define GTM_DUAL__CH0_RX_APT_CFG22A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG22B    32'h00000042
`define GTM_DUAL__CH0_RX_APT_CFG22B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG23A    32'h00000043
`define GTM_DUAL__CH0_RX_APT_CFG23A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG23B    32'h00000044
`define GTM_DUAL__CH0_RX_APT_CFG23B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG24A    32'h00000045
`define GTM_DUAL__CH0_RX_APT_CFG24A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG24B    32'h00000046
`define GTM_DUAL__CH0_RX_APT_CFG24B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG25A    32'h00000047
`define GTM_DUAL__CH0_RX_APT_CFG25A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG25B    32'h00000048
`define GTM_DUAL__CH0_RX_APT_CFG25B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG26A    32'h00000049
`define GTM_DUAL__CH0_RX_APT_CFG26A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG26B    32'h0000004a
`define GTM_DUAL__CH0_RX_APT_CFG26B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG27A    32'h0000004b
`define GTM_DUAL__CH0_RX_APT_CFG27A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG27B    32'h0000004c
`define GTM_DUAL__CH0_RX_APT_CFG27B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG28A    32'h0000004d
`define GTM_DUAL__CH0_RX_APT_CFG28A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG28B    32'h0000004e
`define GTM_DUAL__CH0_RX_APT_CFG28B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG2A    32'h0000004f
`define GTM_DUAL__CH0_RX_APT_CFG2A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG2B    32'h00000050
`define GTM_DUAL__CH0_RX_APT_CFG2B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG3A    32'h00000051
`define GTM_DUAL__CH0_RX_APT_CFG3A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG3B    32'h00000052
`define GTM_DUAL__CH0_RX_APT_CFG3B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG4A    32'h00000053
`define GTM_DUAL__CH0_RX_APT_CFG4A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG4B    32'h00000054
`define GTM_DUAL__CH0_RX_APT_CFG4B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG5A    32'h00000055
`define GTM_DUAL__CH0_RX_APT_CFG5A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG5B    32'h00000056
`define GTM_DUAL__CH0_RX_APT_CFG5B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG6A    32'h00000057
`define GTM_DUAL__CH0_RX_APT_CFG6A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG6B    32'h00000058
`define GTM_DUAL__CH0_RX_APT_CFG6B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG7A    32'h00000059
`define GTM_DUAL__CH0_RX_APT_CFG7A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG7B    32'h0000005a
`define GTM_DUAL__CH0_RX_APT_CFG7B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG8A    32'h0000005b
`define GTM_DUAL__CH0_RX_APT_CFG8A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG8B    32'h0000005c
`define GTM_DUAL__CH0_RX_APT_CFG8B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG9A    32'h0000005d
`define GTM_DUAL__CH0_RX_APT_CFG9A_SZ 16

`define GTM_DUAL__CH0_RX_APT_CFG9B    32'h0000005e
`define GTM_DUAL__CH0_RX_APT_CFG9B_SZ 16

`define GTM_DUAL__CH0_RX_APT_CTRL_CFG2    32'h0000005f
`define GTM_DUAL__CH0_RX_APT_CTRL_CFG2_SZ 16

`define GTM_DUAL__CH0_RX_APT_CTRL_CFG3    32'h00000060
`define GTM_DUAL__CH0_RX_APT_CTRL_CFG3_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG0A    32'h00000061
`define GTM_DUAL__CH0_RX_CAL_CFG0A_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG0B    32'h00000062
`define GTM_DUAL__CH0_RX_CAL_CFG0B_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG1A    32'h00000063
`define GTM_DUAL__CH0_RX_CAL_CFG1A_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG1B    32'h00000064
`define GTM_DUAL__CH0_RX_CAL_CFG1B_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG2A    32'h00000065
`define GTM_DUAL__CH0_RX_CAL_CFG2A_SZ 16

`define GTM_DUAL__CH0_RX_CAL_CFG2B    32'h00000066
`define GTM_DUAL__CH0_RX_CAL_CFG2B_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG0A    32'h00000067
`define GTM_DUAL__CH0_RX_CDR_CFG0A_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG0B    32'h00000068
`define GTM_DUAL__CH0_RX_CDR_CFG0B_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG1A    32'h00000069
`define GTM_DUAL__CH0_RX_CDR_CFG1A_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG1B    32'h0000006a
`define GTM_DUAL__CH0_RX_CDR_CFG1B_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG2A    32'h0000006b
`define GTM_DUAL__CH0_RX_CDR_CFG2A_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG2B    32'h0000006c
`define GTM_DUAL__CH0_RX_CDR_CFG2B_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG3A    32'h0000006d
`define GTM_DUAL__CH0_RX_CDR_CFG3A_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG3B    32'h0000006e
`define GTM_DUAL__CH0_RX_CDR_CFG3B_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG4A    32'h0000006f
`define GTM_DUAL__CH0_RX_CDR_CFG4A_SZ 16

`define GTM_DUAL__CH0_RX_CDR_CFG4B    32'h00000070
`define GTM_DUAL__CH0_RX_CDR_CFG4B_SZ 16

`define GTM_DUAL__CH0_RX_CLKGN_CFG0    32'h00000071
`define GTM_DUAL__CH0_RX_CLKGN_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_CLKGN_CFG1    32'h00000072
`define GTM_DUAL__CH0_RX_CLKGN_CFG1_SZ 16

`define GTM_DUAL__CH0_RX_CTLE_CFG0    32'h00000073
`define GTM_DUAL__CH0_RX_CTLE_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_CTLE_CFG1    32'h00000074
`define GTM_DUAL__CH0_RX_CTLE_CFG1_SZ 16

`define GTM_DUAL__CH0_RX_CTLE_CFG2    32'h00000075
`define GTM_DUAL__CH0_RX_CTLE_CFG2_SZ 16

`define GTM_DUAL__CH0_RX_CTLE_CFG3    32'h00000076
`define GTM_DUAL__CH0_RX_CTLE_CFG3_SZ 16

`define GTM_DUAL__CH0_RX_DSP_CFG    32'h00000077
`define GTM_DUAL__CH0_RX_DSP_CFG_SZ 16

`define GTM_DUAL__CH0_RX_MON_CFG    32'h00000078
`define GTM_DUAL__CH0_RX_MON_CFG_SZ 16

`define GTM_DUAL__CH0_RX_PAD_CFG0    32'h00000079
`define GTM_DUAL__CH0_RX_PAD_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_PAD_CFG1    32'h0000007a
`define GTM_DUAL__CH0_RX_PAD_CFG1_SZ 16

`define GTM_DUAL__CH0_RX_PCS_CFG0    32'h0000007b
`define GTM_DUAL__CH0_RX_PCS_CFG0_SZ 16

`define GTM_DUAL__CH0_RX_PCS_CFG1    32'h0000007c
`define GTM_DUAL__CH0_RX_PCS_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_ANA_CFG0    32'h0000007d
`define GTM_DUAL__CH0_TX_ANA_CFG0_SZ 16

`define GTM_DUAL__CH0_TX_ANA_CFG1    32'h0000007e
`define GTM_DUAL__CH0_TX_ANA_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_ANA_CFG2    32'h0000007f
`define GTM_DUAL__CH0_TX_ANA_CFG2_SZ 16

`define GTM_DUAL__CH0_TX_ANA_CFG3    32'h00000080
`define GTM_DUAL__CH0_TX_ANA_CFG3_SZ 16

`define GTM_DUAL__CH0_TX_ANA_CFG4    32'h00000081
`define GTM_DUAL__CH0_TX_ANA_CFG4_SZ 16

`define GTM_DUAL__CH0_TX_CAL_CFG0    32'h00000082
`define GTM_DUAL__CH0_TX_CAL_CFG0_SZ 16

`define GTM_DUAL__CH0_TX_CAL_CFG1    32'h00000083
`define GTM_DUAL__CH0_TX_CAL_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG0    32'h00000084
`define GTM_DUAL__CH0_TX_DRV_CFG0_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG1    32'h00000085
`define GTM_DUAL__CH0_TX_DRV_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG2    32'h00000086
`define GTM_DUAL__CH0_TX_DRV_CFG2_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG3    32'h00000087
`define GTM_DUAL__CH0_TX_DRV_CFG3_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG4    32'h00000088
`define GTM_DUAL__CH0_TX_DRV_CFG4_SZ 16

`define GTM_DUAL__CH0_TX_DRV_CFG5    32'h00000089
`define GTM_DUAL__CH0_TX_DRV_CFG5_SZ 16

`define GTM_DUAL__CH0_TX_LPBK_CFG0    32'h0000008a
`define GTM_DUAL__CH0_TX_LPBK_CFG0_SZ 16

`define GTM_DUAL__CH0_TX_LPBK_CFG1    32'h0000008b
`define GTM_DUAL__CH0_TX_LPBK_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG0    32'h0000008c
`define GTM_DUAL__CH0_TX_PCS_CFG0_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG1    32'h0000008d
`define GTM_DUAL__CH0_TX_PCS_CFG1_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG10    32'h0000008e
`define GTM_DUAL__CH0_TX_PCS_CFG10_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG11    32'h0000008f
`define GTM_DUAL__CH0_TX_PCS_CFG11_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG12    32'h00000090
`define GTM_DUAL__CH0_TX_PCS_CFG12_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG13    32'h00000091
`define GTM_DUAL__CH0_TX_PCS_CFG13_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG14    32'h00000092
`define GTM_DUAL__CH0_TX_PCS_CFG14_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG15    32'h00000093
`define GTM_DUAL__CH0_TX_PCS_CFG15_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG16    32'h00000094
`define GTM_DUAL__CH0_TX_PCS_CFG16_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG17    32'h00000095
`define GTM_DUAL__CH0_TX_PCS_CFG17_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG2    32'h00000096
`define GTM_DUAL__CH0_TX_PCS_CFG2_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG3    32'h00000097
`define GTM_DUAL__CH0_TX_PCS_CFG3_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG4    32'h00000098
`define GTM_DUAL__CH0_TX_PCS_CFG4_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG5    32'h00000099
`define GTM_DUAL__CH0_TX_PCS_CFG5_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG6    32'h0000009a
`define GTM_DUAL__CH0_TX_PCS_CFG6_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG7    32'h0000009b
`define GTM_DUAL__CH0_TX_PCS_CFG7_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG8    32'h0000009c
`define GTM_DUAL__CH0_TX_PCS_CFG8_SZ 16

`define GTM_DUAL__CH0_TX_PCS_CFG9    32'h0000009d
`define GTM_DUAL__CH0_TX_PCS_CFG9_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG0    32'h0000009e
`define GTM_DUAL__CH1_A_CH_CFG0_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG1    32'h0000009f
`define GTM_DUAL__CH1_A_CH_CFG1_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG2    32'h000000a0
`define GTM_DUAL__CH1_A_CH_CFG2_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG3    32'h000000a1
`define GTM_DUAL__CH1_A_CH_CFG3_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG4    32'h000000a2
`define GTM_DUAL__CH1_A_CH_CFG4_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG5    32'h000000a3
`define GTM_DUAL__CH1_A_CH_CFG5_SZ 16

`define GTM_DUAL__CH1_A_CH_CFG6    32'h000000a4
`define GTM_DUAL__CH1_A_CH_CFG6_SZ 16

`define GTM_DUAL__CH1_RST_LP_CFG0    32'h000000a5
`define GTM_DUAL__CH1_RST_LP_CFG0_SZ 16

`define GTM_DUAL__CH1_RST_LP_CFG1    32'h000000a6
`define GTM_DUAL__CH1_RST_LP_CFG1_SZ 16

`define GTM_DUAL__CH1_RST_LP_CFG2    32'h000000a7
`define GTM_DUAL__CH1_RST_LP_CFG2_SZ 16

`define GTM_DUAL__CH1_RST_LP_CFG3    32'h000000a8
`define GTM_DUAL__CH1_RST_LP_CFG3_SZ 16

`define GTM_DUAL__CH1_RST_LP_CFG4    32'h000000a9
`define GTM_DUAL__CH1_RST_LP_CFG4_SZ 16

`define GTM_DUAL__CH1_RST_LP_ID_CFG0    32'h000000aa
`define GTM_DUAL__CH1_RST_LP_ID_CFG0_SZ 16

`define GTM_DUAL__CH1_RST_LP_ID_CFG1    32'h000000ab
`define GTM_DUAL__CH1_RST_LP_ID_CFG1_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG0    32'h000000ac
`define GTM_DUAL__CH1_RST_TIME_CFG0_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG1    32'h000000ad
`define GTM_DUAL__CH1_RST_TIME_CFG1_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG2    32'h000000ae
`define GTM_DUAL__CH1_RST_TIME_CFG2_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG3    32'h000000af
`define GTM_DUAL__CH1_RST_TIME_CFG3_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG4    32'h000000b0
`define GTM_DUAL__CH1_RST_TIME_CFG4_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG5    32'h000000b1
`define GTM_DUAL__CH1_RST_TIME_CFG5_SZ 16

`define GTM_DUAL__CH1_RST_TIME_CFG6    32'h000000b2
`define GTM_DUAL__CH1_RST_TIME_CFG6_SZ 16

`define GTM_DUAL__CH1_RX_ADC_CFG0    32'h000000b3
`define GTM_DUAL__CH1_RX_ADC_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_ADC_CFG1    32'h000000b4
`define GTM_DUAL__CH1_RX_ADC_CFG1_SZ 16

`define GTM_DUAL__CH1_RX_ANA_CFG0    32'h000000b5
`define GTM_DUAL__CH1_RX_ANA_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_ANA_CFG1    32'h000000b6
`define GTM_DUAL__CH1_RX_ANA_CFG1_SZ 16

`define GTM_DUAL__CH1_RX_ANA_CFG2    32'h000000b7
`define GTM_DUAL__CH1_RX_ANA_CFG2_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG0A    32'h000000b8
`define GTM_DUAL__CH1_RX_APT_CFG0A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG0B    32'h000000b9
`define GTM_DUAL__CH1_RX_APT_CFG0B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG10A    32'h000000ba
`define GTM_DUAL__CH1_RX_APT_CFG10A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG10B    32'h000000bb
`define GTM_DUAL__CH1_RX_APT_CFG10B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG11A    32'h000000bc
`define GTM_DUAL__CH1_RX_APT_CFG11A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG11B    32'h000000bd
`define GTM_DUAL__CH1_RX_APT_CFG11B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG12A    32'h000000be
`define GTM_DUAL__CH1_RX_APT_CFG12A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG12B    32'h000000bf
`define GTM_DUAL__CH1_RX_APT_CFG12B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG13A    32'h000000c0
`define GTM_DUAL__CH1_RX_APT_CFG13A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG13B    32'h000000c1
`define GTM_DUAL__CH1_RX_APT_CFG13B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG14A    32'h000000c2
`define GTM_DUAL__CH1_RX_APT_CFG14A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG14B    32'h000000c3
`define GTM_DUAL__CH1_RX_APT_CFG14B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG15A    32'h000000c4
`define GTM_DUAL__CH1_RX_APT_CFG15A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG15B    32'h000000c5
`define GTM_DUAL__CH1_RX_APT_CFG15B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG16A    32'h000000c6
`define GTM_DUAL__CH1_RX_APT_CFG16A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG16B    32'h000000c7
`define GTM_DUAL__CH1_RX_APT_CFG16B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG17A    32'h000000c8
`define GTM_DUAL__CH1_RX_APT_CFG17A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG17B    32'h000000c9
`define GTM_DUAL__CH1_RX_APT_CFG17B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG18A    32'h000000ca
`define GTM_DUAL__CH1_RX_APT_CFG18A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG18B    32'h000000cb
`define GTM_DUAL__CH1_RX_APT_CFG18B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG19A    32'h000000cc
`define GTM_DUAL__CH1_RX_APT_CFG19A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG19B    32'h000000cd
`define GTM_DUAL__CH1_RX_APT_CFG19B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG1A    32'h000000ce
`define GTM_DUAL__CH1_RX_APT_CFG1A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG1B    32'h000000cf
`define GTM_DUAL__CH1_RX_APT_CFG1B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG20A    32'h000000d0
`define GTM_DUAL__CH1_RX_APT_CFG20A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG20B    32'h000000d1
`define GTM_DUAL__CH1_RX_APT_CFG20B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG21A    32'h000000d2
`define GTM_DUAL__CH1_RX_APT_CFG21A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG21B    32'h000000d3
`define GTM_DUAL__CH1_RX_APT_CFG21B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG22A    32'h000000d4
`define GTM_DUAL__CH1_RX_APT_CFG22A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG22B    32'h000000d5
`define GTM_DUAL__CH1_RX_APT_CFG22B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG23A    32'h000000d6
`define GTM_DUAL__CH1_RX_APT_CFG23A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG23B    32'h000000d7
`define GTM_DUAL__CH1_RX_APT_CFG23B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG24A    32'h000000d8
`define GTM_DUAL__CH1_RX_APT_CFG24A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG24B    32'h000000d9
`define GTM_DUAL__CH1_RX_APT_CFG24B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG25A    32'h000000da
`define GTM_DUAL__CH1_RX_APT_CFG25A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG25B    32'h000000db
`define GTM_DUAL__CH1_RX_APT_CFG25B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG26A    32'h000000dc
`define GTM_DUAL__CH1_RX_APT_CFG26A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG26B    32'h000000dd
`define GTM_DUAL__CH1_RX_APT_CFG26B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG27A    32'h000000de
`define GTM_DUAL__CH1_RX_APT_CFG27A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG27B    32'h000000df
`define GTM_DUAL__CH1_RX_APT_CFG27B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG28A    32'h000000e0
`define GTM_DUAL__CH1_RX_APT_CFG28A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG28B    32'h000000e1
`define GTM_DUAL__CH1_RX_APT_CFG28B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG2A    32'h000000e2
`define GTM_DUAL__CH1_RX_APT_CFG2A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG2B    32'h000000e3
`define GTM_DUAL__CH1_RX_APT_CFG2B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG3A    32'h000000e4
`define GTM_DUAL__CH1_RX_APT_CFG3A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG3B    32'h000000e5
`define GTM_DUAL__CH1_RX_APT_CFG3B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG4A    32'h000000e6
`define GTM_DUAL__CH1_RX_APT_CFG4A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG4B    32'h000000e7
`define GTM_DUAL__CH1_RX_APT_CFG4B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG5A    32'h000000e8
`define GTM_DUAL__CH1_RX_APT_CFG5A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG5B    32'h000000e9
`define GTM_DUAL__CH1_RX_APT_CFG5B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG6A    32'h000000ea
`define GTM_DUAL__CH1_RX_APT_CFG6A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG6B    32'h000000eb
`define GTM_DUAL__CH1_RX_APT_CFG6B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG7A    32'h000000ec
`define GTM_DUAL__CH1_RX_APT_CFG7A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG7B    32'h000000ed
`define GTM_DUAL__CH1_RX_APT_CFG7B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG8A    32'h000000ee
`define GTM_DUAL__CH1_RX_APT_CFG8A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG8B    32'h000000ef
`define GTM_DUAL__CH1_RX_APT_CFG8B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG9A    32'h000000f0
`define GTM_DUAL__CH1_RX_APT_CFG9A_SZ 16

`define GTM_DUAL__CH1_RX_APT_CFG9B    32'h000000f1
`define GTM_DUAL__CH1_RX_APT_CFG9B_SZ 16

`define GTM_DUAL__CH1_RX_APT_CTRL_CFG2    32'h000000f2
`define GTM_DUAL__CH1_RX_APT_CTRL_CFG2_SZ 16

`define GTM_DUAL__CH1_RX_APT_CTRL_CFG3    32'h000000f3
`define GTM_DUAL__CH1_RX_APT_CTRL_CFG3_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG0A    32'h000000f4
`define GTM_DUAL__CH1_RX_CAL_CFG0A_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG0B    32'h000000f5
`define GTM_DUAL__CH1_RX_CAL_CFG0B_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG1A    32'h000000f6
`define GTM_DUAL__CH1_RX_CAL_CFG1A_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG1B    32'h000000f7
`define GTM_DUAL__CH1_RX_CAL_CFG1B_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG2A    32'h000000f8
`define GTM_DUAL__CH1_RX_CAL_CFG2A_SZ 16

`define GTM_DUAL__CH1_RX_CAL_CFG2B    32'h000000f9
`define GTM_DUAL__CH1_RX_CAL_CFG2B_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG0A    32'h000000fa
`define GTM_DUAL__CH1_RX_CDR_CFG0A_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG0B    32'h000000fb
`define GTM_DUAL__CH1_RX_CDR_CFG0B_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG1A    32'h000000fc
`define GTM_DUAL__CH1_RX_CDR_CFG1A_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG1B    32'h000000fd
`define GTM_DUAL__CH1_RX_CDR_CFG1B_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG2A    32'h000000fe
`define GTM_DUAL__CH1_RX_CDR_CFG2A_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG2B    32'h000000ff
`define GTM_DUAL__CH1_RX_CDR_CFG2B_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG3A    32'h00000100
`define GTM_DUAL__CH1_RX_CDR_CFG3A_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG3B    32'h00000101
`define GTM_DUAL__CH1_RX_CDR_CFG3B_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG4A    32'h00000102
`define GTM_DUAL__CH1_RX_CDR_CFG4A_SZ 16

`define GTM_DUAL__CH1_RX_CDR_CFG4B    32'h00000103
`define GTM_DUAL__CH1_RX_CDR_CFG4B_SZ 16

`define GTM_DUAL__CH1_RX_CLKGN_CFG0    32'h00000104
`define GTM_DUAL__CH1_RX_CLKGN_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_CLKGN_CFG1    32'h00000105
`define GTM_DUAL__CH1_RX_CLKGN_CFG1_SZ 16

`define GTM_DUAL__CH1_RX_CTLE_CFG0    32'h00000106
`define GTM_DUAL__CH1_RX_CTLE_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_CTLE_CFG1    32'h00000107
`define GTM_DUAL__CH1_RX_CTLE_CFG1_SZ 16

`define GTM_DUAL__CH1_RX_CTLE_CFG2    32'h00000108
`define GTM_DUAL__CH1_RX_CTLE_CFG2_SZ 16

`define GTM_DUAL__CH1_RX_CTLE_CFG3    32'h00000109
`define GTM_DUAL__CH1_RX_CTLE_CFG3_SZ 16

`define GTM_DUAL__CH1_RX_DSP_CFG    32'h0000010a
`define GTM_DUAL__CH1_RX_DSP_CFG_SZ 16

`define GTM_DUAL__CH1_RX_MON_CFG    32'h0000010b
`define GTM_DUAL__CH1_RX_MON_CFG_SZ 16

`define GTM_DUAL__CH1_RX_PAD_CFG0    32'h0000010c
`define GTM_DUAL__CH1_RX_PAD_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_PAD_CFG1    32'h0000010d
`define GTM_DUAL__CH1_RX_PAD_CFG1_SZ 16

`define GTM_DUAL__CH1_RX_PCS_CFG0    32'h0000010e
`define GTM_DUAL__CH1_RX_PCS_CFG0_SZ 16

`define GTM_DUAL__CH1_RX_PCS_CFG1    32'h0000010f
`define GTM_DUAL__CH1_RX_PCS_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_ANA_CFG0    32'h00000110
`define GTM_DUAL__CH1_TX_ANA_CFG0_SZ 16

`define GTM_DUAL__CH1_TX_ANA_CFG1    32'h00000111
`define GTM_DUAL__CH1_TX_ANA_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_ANA_CFG2    32'h00000112
`define GTM_DUAL__CH1_TX_ANA_CFG2_SZ 16

`define GTM_DUAL__CH1_TX_ANA_CFG3    32'h00000113
`define GTM_DUAL__CH1_TX_ANA_CFG3_SZ 16

`define GTM_DUAL__CH1_TX_ANA_CFG4    32'h00000114
`define GTM_DUAL__CH1_TX_ANA_CFG4_SZ 16

`define GTM_DUAL__CH1_TX_CAL_CFG0    32'h00000115
`define GTM_DUAL__CH1_TX_CAL_CFG0_SZ 16

`define GTM_DUAL__CH1_TX_CAL_CFG1    32'h00000116
`define GTM_DUAL__CH1_TX_CAL_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG0    32'h00000117
`define GTM_DUAL__CH1_TX_DRV_CFG0_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG1    32'h00000118
`define GTM_DUAL__CH1_TX_DRV_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG2    32'h00000119
`define GTM_DUAL__CH1_TX_DRV_CFG2_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG3    32'h0000011a
`define GTM_DUAL__CH1_TX_DRV_CFG3_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG4    32'h0000011b
`define GTM_DUAL__CH1_TX_DRV_CFG4_SZ 16

`define GTM_DUAL__CH1_TX_DRV_CFG5    32'h0000011c
`define GTM_DUAL__CH1_TX_DRV_CFG5_SZ 16

`define GTM_DUAL__CH1_TX_LPBK_CFG0    32'h0000011d
`define GTM_DUAL__CH1_TX_LPBK_CFG0_SZ 16

`define GTM_DUAL__CH1_TX_LPBK_CFG1    32'h0000011e
`define GTM_DUAL__CH1_TX_LPBK_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG0    32'h0000011f
`define GTM_DUAL__CH1_TX_PCS_CFG0_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG1    32'h00000120
`define GTM_DUAL__CH1_TX_PCS_CFG1_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG10    32'h00000121
`define GTM_DUAL__CH1_TX_PCS_CFG10_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG11    32'h00000122
`define GTM_DUAL__CH1_TX_PCS_CFG11_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG12    32'h00000123
`define GTM_DUAL__CH1_TX_PCS_CFG12_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG13    32'h00000124
`define GTM_DUAL__CH1_TX_PCS_CFG13_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG14    32'h00000125
`define GTM_DUAL__CH1_TX_PCS_CFG14_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG15    32'h00000126
`define GTM_DUAL__CH1_TX_PCS_CFG15_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG16    32'h00000127
`define GTM_DUAL__CH1_TX_PCS_CFG16_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG17    32'h00000128
`define GTM_DUAL__CH1_TX_PCS_CFG17_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG2    32'h00000129
`define GTM_DUAL__CH1_TX_PCS_CFG2_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG3    32'h0000012a
`define GTM_DUAL__CH1_TX_PCS_CFG3_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG4    32'h0000012b
`define GTM_DUAL__CH1_TX_PCS_CFG4_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG5    32'h0000012c
`define GTM_DUAL__CH1_TX_PCS_CFG5_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG6    32'h0000012d
`define GTM_DUAL__CH1_TX_PCS_CFG6_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG7    32'h0000012e
`define GTM_DUAL__CH1_TX_PCS_CFG7_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG8    32'h0000012f
`define GTM_DUAL__CH1_TX_PCS_CFG8_SZ 16

`define GTM_DUAL__CH1_TX_PCS_CFG9    32'h00000130
`define GTM_DUAL__CH1_TX_PCS_CFG9_SZ 16

`define GTM_DUAL__DATARATE    32'h00000131
`define GTM_DUAL__DATARATE_SZ 64

`define GTM_DUAL__DRPEN_CFG    32'h00000132
`define GTM_DUAL__DRPEN_CFG_SZ 16

`define GTM_DUAL__FEC_CFG0    32'h00000133
`define GTM_DUAL__FEC_CFG0_SZ 16

`define GTM_DUAL__FEC_CFG1    32'h00000134
`define GTM_DUAL__FEC_CFG1_SZ 16

`define GTM_DUAL__FEC_CFG10    32'h00000135
`define GTM_DUAL__FEC_CFG10_SZ 16

`define GTM_DUAL__FEC_CFG11    32'h00000136
`define GTM_DUAL__FEC_CFG11_SZ 16

`define GTM_DUAL__FEC_CFG12    32'h00000137
`define GTM_DUAL__FEC_CFG12_SZ 16

`define GTM_DUAL__FEC_CFG13    32'h00000138
`define GTM_DUAL__FEC_CFG13_SZ 16

`define GTM_DUAL__FEC_CFG14    32'h00000139
`define GTM_DUAL__FEC_CFG14_SZ 16

`define GTM_DUAL__FEC_CFG15    32'h0000013a
`define GTM_DUAL__FEC_CFG15_SZ 16

`define GTM_DUAL__FEC_CFG16    32'h0000013b
`define GTM_DUAL__FEC_CFG16_SZ 16

`define GTM_DUAL__FEC_CFG17    32'h0000013c
`define GTM_DUAL__FEC_CFG17_SZ 16

`define GTM_DUAL__FEC_CFG18    32'h0000013d
`define GTM_DUAL__FEC_CFG18_SZ 16

`define GTM_DUAL__FEC_CFG19    32'h0000013e
`define GTM_DUAL__FEC_CFG19_SZ 16

`define GTM_DUAL__FEC_CFG2    32'h0000013f
`define GTM_DUAL__FEC_CFG2_SZ 16

`define GTM_DUAL__FEC_CFG20    32'h00000140
`define GTM_DUAL__FEC_CFG20_SZ 16

`define GTM_DUAL__FEC_CFG21    32'h00000141
`define GTM_DUAL__FEC_CFG21_SZ 16

`define GTM_DUAL__FEC_CFG22    32'h00000142
`define GTM_DUAL__FEC_CFG22_SZ 16

`define GTM_DUAL__FEC_CFG23    32'h00000143
`define GTM_DUAL__FEC_CFG23_SZ 16

`define GTM_DUAL__FEC_CFG24    32'h00000144
`define GTM_DUAL__FEC_CFG24_SZ 16

`define GTM_DUAL__FEC_CFG25    32'h00000145
`define GTM_DUAL__FEC_CFG25_SZ 16

`define GTM_DUAL__FEC_CFG26    32'h00000146
`define GTM_DUAL__FEC_CFG26_SZ 16

`define GTM_DUAL__FEC_CFG27    32'h00000147
`define GTM_DUAL__FEC_CFG27_SZ 16

`define GTM_DUAL__FEC_CFG3    32'h00000148
`define GTM_DUAL__FEC_CFG3_SZ 16

`define GTM_DUAL__FEC_CFG4    32'h00000149
`define GTM_DUAL__FEC_CFG4_SZ 16

`define GTM_DUAL__FEC_CFG5    32'h0000014a
`define GTM_DUAL__FEC_CFG5_SZ 16

`define GTM_DUAL__FEC_CFG6    32'h0000014b
`define GTM_DUAL__FEC_CFG6_SZ 16

`define GTM_DUAL__FEC_CFG7    32'h0000014c
`define GTM_DUAL__FEC_CFG7_SZ 16

`define GTM_DUAL__FEC_CFG8    32'h0000014d
`define GTM_DUAL__FEC_CFG8_SZ 16

`define GTM_DUAL__FEC_CFG9    32'h0000014e
`define GTM_DUAL__FEC_CFG9_SZ 16

`define GTM_DUAL__FEC_MODE    32'h0000014f
`define GTM_DUAL__FEC_MODE_SZ 48

`define GTM_DUAL__INS_LOSS_NYQ    32'h00000150
`define GTM_DUAL__INS_LOSS_NYQ_SZ 64

`define GTM_DUAL__INTERFACE_WIDTH    32'h00000151
`define GTM_DUAL__INTERFACE_WIDTH_SZ 9

`define GTM_DUAL__MODULATION_MODE    32'h00000152
`define GTM_DUAL__MODULATION_MODE_SZ 32

`define GTM_DUAL__PLL_CFG0    32'h00000153
`define GTM_DUAL__PLL_CFG0_SZ 16

`define GTM_DUAL__PLL_CFG1    32'h00000154
`define GTM_DUAL__PLL_CFG1_SZ 16

`define GTM_DUAL__PLL_CFG2    32'h00000155
`define GTM_DUAL__PLL_CFG2_SZ 16

`define GTM_DUAL__PLL_CFG3    32'h00000156
`define GTM_DUAL__PLL_CFG3_SZ 16

`define GTM_DUAL__PLL_CFG4    32'h00000157
`define GTM_DUAL__PLL_CFG4_SZ 16

`define GTM_DUAL__PLL_CFG5    32'h00000158
`define GTM_DUAL__PLL_CFG5_SZ 16

`define GTM_DUAL__PLL_CFG6    32'h00000159
`define GTM_DUAL__PLL_CFG6_SZ 16

`define GTM_DUAL__PLL_CRS_CTRL_CFG0    32'h0000015a
`define GTM_DUAL__PLL_CRS_CTRL_CFG0_SZ 16

`define GTM_DUAL__PLL_CRS_CTRL_CFG1    32'h0000015b
`define GTM_DUAL__PLL_CRS_CTRL_CFG1_SZ 16

`define GTM_DUAL__PLL_IPS_PIN_EN    32'h0000015c
`define GTM_DUAL__PLL_IPS_PIN_EN_SZ 1

`define GTM_DUAL__PLL_IPS_REFCLK_SEL    32'h0000015d
`define GTM_DUAL__PLL_IPS_REFCLK_SEL_SZ 3

`define GTM_DUAL__RCALSAP_TESTEN    32'h0000015e
`define GTM_DUAL__RCALSAP_TESTEN_SZ 1

`define GTM_DUAL__RCAL_APROBE    32'h0000015f
`define GTM_DUAL__RCAL_APROBE_SZ 1

`define GTM_DUAL__RST_CFG    32'h00000160
`define GTM_DUAL__RST_CFG_SZ 16

`define GTM_DUAL__RST_PLL_CFG0    32'h00000161
`define GTM_DUAL__RST_PLL_CFG0_SZ 16

`define GTM_DUAL__SAP_CFG0    32'h00000162
`define GTM_DUAL__SAP_CFG0_SZ 16

`define GTM_DUAL__SDM_CFG0    32'h00000163
`define GTM_DUAL__SDM_CFG0_SZ 16

`define GTM_DUAL__SDM_CFG1    32'h00000164
`define GTM_DUAL__SDM_CFG1_SZ 16

`define GTM_DUAL__SDM_CFG2    32'h00000165
`define GTM_DUAL__SDM_CFG2_SZ 16

`define GTM_DUAL__SDM_SEED_CFG0    32'h00000166
`define GTM_DUAL__SDM_SEED_CFG0_SZ 16

`define GTM_DUAL__SDM_SEED_CFG1    32'h00000167
`define GTM_DUAL__SDM_SEED_CFG1_SZ 16

`define GTM_DUAL__SIM_DEVICE    32'h00000168
`define GTM_DUAL__SIM_DEVICE_SZ 152

`define GTM_DUAL__SIM_RESET_SPEEDUP    32'h00000169
`define GTM_DUAL__SIM_RESET_SPEEDUP_SZ 40

`define GTM_DUAL__TX_AMPLITUDE_SWING    32'h0000016a
`define GTM_DUAL__TX_AMPLITUDE_SWING_SZ 11

`endif  // B_GTM_DUAL_DEFINES_VH