// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HNICPIPE_QUAD_DEFINES_VH
`else
`define B_HNICPIPE_QUAD_DEFINES_VH

// Look-up table parameters
//

`define HNICPIPE_QUAD_ADDR_N  16
`define HNICPIPE_QUAD_ADDR_SZ 32
`define HNICPIPE_QUAD_DATA_SZ 32

// Attribute addresses
//

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG0    32'h00000000
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG0_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG1    32'h00000001
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG1_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG2    32'h00000002
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG2_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG3    32'h00000003
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG3_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG4    32'h00000004
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG4_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG5    32'h00000005
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG5_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG6    32'h00000006
`define HNICPIPE_QUAD__HNICPIPE_HPIPE_CFG6_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_OPTDLY_CFG0    32'h00000007
`define HNICPIPE_QUAD__HNICPIPE_OPTDLY_CFG0_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_OPTDLY_CFG1    32'h00000008
`define HNICPIPE_QUAD__HNICPIPE_OPTDLY_CFG1_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_PIPE_CFG    32'h00000009
`define HNICPIPE_QUAD__HNICPIPE_PIPE_CFG_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_RX_CLKMUX_SEL    32'h0000000a
`define HNICPIPE_QUAD__HNICPIPE_RX_CLKMUX_SEL_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_RX_CLK_REMAP_CFG    32'h0000000b
`define HNICPIPE_QUAD__HNICPIPE_RX_CLK_REMAP_CFG_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_RX_DATA_REMAP_CFG    32'h0000000c
`define HNICPIPE_QUAD__HNICPIPE_RX_DATA_REMAP_CFG_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_TX_CLKMUX_SEL    32'h0000000d
`define HNICPIPE_QUAD__HNICPIPE_TX_CLKMUX_SEL_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_TX_CLK_REMAP_CFG    32'h0000000e
`define HNICPIPE_QUAD__HNICPIPE_TX_CLK_REMAP_CFG_SZ 32

`define HNICPIPE_QUAD__HNICPIPE_TX_DATA_REMAP_CFG    32'h0000000f
`define HNICPIPE_QUAD__HNICPIPE_TX_DATA_REMAP_CFG_SZ 32

`endif  // B_HNICPIPE_QUAD_DEFINES_VH