`include "B_IDELAYE2_defines.vh"

reg [`IDELAYE2_DATA_SZ-1:0] ATTR [0:`IDELAYE2_ADDR_N-1];
reg [`IDELAYE2__CINVCTRL_SEL_SZ:1] CINVCTRL_SEL_REG = CINVCTRL_SEL;
reg [`IDELAYE2__DELAY_SRC_SZ:1] DELAY_SRC_REG = DELAY_SRC;
reg [`IDELAYE2__HIGH_PERFORMANCE_MODE_SZ:1] HIGH_PERFORMANCE_MODE_REG = HIGH_PERFORMANCE_MODE;
reg [`IDELAYE2__IDELAY_TYPE_SZ:1] IDELAY_TYPE_REG = IDELAY_TYPE;
reg [`IDELAYE2__IDELAY_VALUE_SZ-1:0] IDELAY_VALUE_REG = IDELAY_VALUE;
reg IS_C_INVERTED_REG = IS_C_INVERTED;
reg IS_DATAIN_INVERTED_REG = IS_DATAIN_INVERTED;
reg IS_IDATAIN_INVERTED_REG = IS_IDATAIN_INVERTED;
reg [`IDELAYE2__PIPE_SEL_SZ:1] PIPE_SEL_REG = PIPE_SEL;
real REFCLK_FREQUENCY_REG = REFCLK_FREQUENCY;
reg [`IDELAYE2__SIGNAL_PATTERN_SZ:1] SIGNAL_PATTERN_REG = SIGNAL_PATTERN;
reg [`IDELAYE2__SIM_DELAY_D_SZ-1:0] SIM_DELAY_D_REG = SIM_DELAY_D;

initial begin
  ATTR[`IDELAYE2__CINVCTRL_SEL] = CINVCTRL_SEL;
  ATTR[`IDELAYE2__DELAY_SRC] = DELAY_SRC;
  ATTR[`IDELAYE2__HIGH_PERFORMANCE_MODE] = HIGH_PERFORMANCE_MODE;
  ATTR[`IDELAYE2__IDELAY_TYPE] = IDELAY_TYPE;
  ATTR[`IDELAYE2__IDELAY_VALUE] = IDELAY_VALUE;
  ATTR[`IDELAYE2__IS_C_INVERTED] = IS_C_INVERTED;
  ATTR[`IDELAYE2__IS_DATAIN_INVERTED] = IS_DATAIN_INVERTED;
  ATTR[`IDELAYE2__IS_IDATAIN_INVERTED] = IS_IDATAIN_INVERTED;
  ATTR[`IDELAYE2__PIPE_SEL] = PIPE_SEL;
  ATTR[`IDELAYE2__REFCLK_FREQUENCY] = $realtobits(REFCLK_FREQUENCY);
  ATTR[`IDELAYE2__SIGNAL_PATTERN] = SIGNAL_PATTERN;
  ATTR[`IDELAYE2__SIM_DELAY_D] = SIM_DELAY_D;
end

always @(trig_attr) begin
  CINVCTRL_SEL_REG = ATTR[`IDELAYE2__CINVCTRL_SEL];
  DELAY_SRC_REG = ATTR[`IDELAYE2__DELAY_SRC];
  HIGH_PERFORMANCE_MODE_REG = ATTR[`IDELAYE2__HIGH_PERFORMANCE_MODE];
  IDELAY_TYPE_REG = ATTR[`IDELAYE2__IDELAY_TYPE];
  IDELAY_VALUE_REG = ATTR[`IDELAYE2__IDELAY_VALUE];
  IS_C_INVERTED_REG = ATTR[`IDELAYE2__IS_C_INVERTED];
  IS_DATAIN_INVERTED_REG = ATTR[`IDELAYE2__IS_DATAIN_INVERTED];
  IS_IDATAIN_INVERTED_REG = ATTR[`IDELAYE2__IS_IDATAIN_INVERTED];
  PIPE_SEL_REG = ATTR[`IDELAYE2__PIPE_SEL];
  REFCLK_FREQUENCY_REG = $bitstoreal(ATTR[`IDELAYE2__REFCLK_FREQUENCY]);
  SIGNAL_PATTERN_REG = ATTR[`IDELAYE2__SIGNAL_PATTERN];
  SIM_DELAY_D_REG = ATTR[`IDELAYE2__SIM_DELAY_D];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IDELAYE2_ADDR_SZ-1:0] addr;
  input  [`IDELAYE2_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IDELAYE2_DATA_SZ-1:0] read_attr;
  input  [`IDELAYE2_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
