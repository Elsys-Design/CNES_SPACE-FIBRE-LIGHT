// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_XPHY_DEFINES_VH
`else
`define B_XPHY_DEFINES_VH

// Look-up table parameters
//

`define XPHY_ADDR_N  88
`define XPHY_ADDR_SZ 32
`define XPHY_DATA_SZ 104

// Attribute addresses
//

`define XPHY__CASCADE_0    32'h00000000
`define XPHY__CASCADE_0_SZ 40

`define XPHY__CASCADE_1    32'h00000001
`define XPHY__CASCADE_1_SZ 40

`define XPHY__CASCADE_2    32'h00000002
`define XPHY__CASCADE_2_SZ 40

`define XPHY__CASCADE_3    32'h00000003
`define XPHY__CASCADE_3_SZ 40

`define XPHY__CASCADE_4    32'h00000004
`define XPHY__CASCADE_4_SZ 40

`define XPHY__CASCADE_5    32'h00000005
`define XPHY__CASCADE_5_SZ 40

`define XPHY__CONTINUOUS_DQS    32'h00000006
`define XPHY__CONTINUOUS_DQS_SZ 40

`define XPHY__CRSE_DLY_EN    32'h00000007
`define XPHY__CRSE_DLY_EN_SZ 40

`define XPHY__DELAY_VALUE_0    32'h00000008
`define XPHY__DELAY_VALUE_0_SZ 11

`define XPHY__DELAY_VALUE_1    32'h00000009
`define XPHY__DELAY_VALUE_1_SZ 11

`define XPHY__DELAY_VALUE_2    32'h0000000a
`define XPHY__DELAY_VALUE_2_SZ 11

`define XPHY__DELAY_VALUE_3    32'h0000000b
`define XPHY__DELAY_VALUE_3_SZ 11

`define XPHY__DELAY_VALUE_4    32'h0000000c
`define XPHY__DELAY_VALUE_4_SZ 11

`define XPHY__DELAY_VALUE_5    32'h0000000d
`define XPHY__DELAY_VALUE_5_SZ 11

`define XPHY__DIS_IDLY_VT_TRACK    32'h0000000e
`define XPHY__DIS_IDLY_VT_TRACK_SZ 40

`define XPHY__DIS_ODLY_VT_TRACK    32'h0000000f
`define XPHY__DIS_ODLY_VT_TRACK_SZ 40

`define XPHY__DIS_QDLY_VT_TRACK    32'h00000010
`define XPHY__DIS_QDLY_VT_TRACK_SZ 40

`define XPHY__DQS_MODE    32'h00000011
`define XPHY__DQS_MODE_SZ 104

`define XPHY__DQS_SRC    32'h00000012
`define XPHY__DQS_SRC_SZ 48

`define XPHY__EN_CLK_TO_LOWER    32'h00000013
`define XPHY__EN_CLK_TO_LOWER_SZ 56

`define XPHY__EN_CLK_TO_UPPER    32'h00000014
`define XPHY__EN_CLK_TO_UPPER_SZ 56

`define XPHY__EN_DYN_DLY_MODE    32'h00000015
`define XPHY__EN_DYN_DLY_MODE_SZ 40

`define XPHY__EN_OTHER_NCLK    32'h00000016
`define XPHY__EN_OTHER_NCLK_SZ 40

`define XPHY__EN_OTHER_PCLK    32'h00000017
`define XPHY__EN_OTHER_PCLK_SZ 40

`define XPHY__FAST_CK    32'h00000018
`define XPHY__FAST_CK_SZ 40

`define XPHY__FIFO_MODE_0    32'h00000019
`define XPHY__FIFO_MODE_0_SZ 48

`define XPHY__FIFO_MODE_1    32'h0000001a
`define XPHY__FIFO_MODE_1_SZ 48

`define XPHY__FIFO_MODE_2    32'h0000001b
`define XPHY__FIFO_MODE_2_SZ 48

`define XPHY__FIFO_MODE_3    32'h0000001c
`define XPHY__FIFO_MODE_3_SZ 48

`define XPHY__FIFO_MODE_4    32'h0000001d
`define XPHY__FIFO_MODE_4_SZ 48

`define XPHY__FIFO_MODE_5    32'h0000001e
`define XPHY__FIFO_MODE_5_SZ 48

`define XPHY__IBUF_DIS_SRC_0    32'h0000001f
`define XPHY__IBUF_DIS_SRC_0_SZ 64

`define XPHY__IBUF_DIS_SRC_1    32'h00000020
`define XPHY__IBUF_DIS_SRC_1_SZ 64

`define XPHY__IBUF_DIS_SRC_2    32'h00000021
`define XPHY__IBUF_DIS_SRC_2_SZ 64

`define XPHY__IBUF_DIS_SRC_3    32'h00000022
`define XPHY__IBUF_DIS_SRC_3_SZ 64

`define XPHY__IBUF_DIS_SRC_4    32'h00000023
`define XPHY__IBUF_DIS_SRC_4_SZ 64

`define XPHY__IBUF_DIS_SRC_5    32'h00000024
`define XPHY__IBUF_DIS_SRC_5_SZ 64

`define XPHY__INV_RXCLK    32'h00000025
`define XPHY__INV_RXCLK_SZ 40

`define XPHY__LP4_DQS    32'h00000026
`define XPHY__LP4_DQS_SZ 40

`define XPHY__ODELAY_BYPASS_0    32'h00000027
`define XPHY__ODELAY_BYPASS_0_SZ 40

`define XPHY__ODELAY_BYPASS_1    32'h00000028
`define XPHY__ODELAY_BYPASS_1_SZ 40

`define XPHY__ODELAY_BYPASS_2    32'h00000029
`define XPHY__ODELAY_BYPASS_2_SZ 40

`define XPHY__ODELAY_BYPASS_3    32'h0000002a
`define XPHY__ODELAY_BYPASS_3_SZ 40

`define XPHY__ODELAY_BYPASS_4    32'h0000002b
`define XPHY__ODELAY_BYPASS_4_SZ 40

`define XPHY__ODELAY_BYPASS_5    32'h0000002c
`define XPHY__ODELAY_BYPASS_5_SZ 40

`define XPHY__ODT_SRC_0    32'h0000002d
`define XPHY__ODT_SRC_0_SZ 64

`define XPHY__ODT_SRC_1    32'h0000002e
`define XPHY__ODT_SRC_1_SZ 64

`define XPHY__ODT_SRC_2    32'h0000002f
`define XPHY__ODT_SRC_2_SZ 64

`define XPHY__ODT_SRC_3    32'h00000030
`define XPHY__ODT_SRC_3_SZ 64

`define XPHY__ODT_SRC_4    32'h00000031
`define XPHY__ODT_SRC_4_SZ 64

`define XPHY__ODT_SRC_5    32'h00000032
`define XPHY__ODT_SRC_5_SZ 64

`define XPHY__PRIME_VAL    32'h00000033
`define XPHY__PRIME_VAL_SZ 1

`define XPHY__REFCLK_FREQUENCY    32'h00000034
`define XPHY__REFCLK_FREQUENCY_SZ 64

`define XPHY__RX_CLK_PHASE_N    32'h00000035
`define XPHY__RX_CLK_PHASE_N_SZ 64

`define XPHY__RX_CLK_PHASE_P    32'h00000036
`define XPHY__RX_CLK_PHASE_P_SZ 64

`define XPHY__RX_DATA_WIDTH    32'h00000037
`define XPHY__RX_DATA_WIDTH_SZ 4

`define XPHY__RX_GATING    32'h00000038
`define XPHY__RX_GATING_SZ 56

`define XPHY__SELF_CALIBRATE    32'h00000039
`define XPHY__SELF_CALIBRATE_SZ 56

`define XPHY__SERIAL_MODE    32'h0000003a
`define XPHY__SERIAL_MODE_SZ 40

`define XPHY__TBYTE_CTL_0    32'h0000003b
`define XPHY__TBYTE_CTL_0_SZ 64

`define XPHY__TBYTE_CTL_1    32'h0000003c
`define XPHY__TBYTE_CTL_1_SZ 64

`define XPHY__TBYTE_CTL_2    32'h0000003d
`define XPHY__TBYTE_CTL_2_SZ 64

`define XPHY__TBYTE_CTL_3    32'h0000003e
`define XPHY__TBYTE_CTL_3_SZ 64

`define XPHY__TBYTE_CTL_4    32'h0000003f
`define XPHY__TBYTE_CTL_4_SZ 64

`define XPHY__TBYTE_CTL_5    32'h00000040
`define XPHY__TBYTE_CTL_5_SZ 64

`define XPHY__TXRX_LOOPBACK_0    32'h00000041
`define XPHY__TXRX_LOOPBACK_0_SZ 40

`define XPHY__TXRX_LOOPBACK_1    32'h00000042
`define XPHY__TXRX_LOOPBACK_1_SZ 40

`define XPHY__TXRX_LOOPBACK_2    32'h00000043
`define XPHY__TXRX_LOOPBACK_2_SZ 40

`define XPHY__TXRX_LOOPBACK_3    32'h00000044
`define XPHY__TXRX_LOOPBACK_3_SZ 40

`define XPHY__TXRX_LOOPBACK_4    32'h00000045
`define XPHY__TXRX_LOOPBACK_4_SZ 40

`define XPHY__TXRX_LOOPBACK_5    32'h00000046
`define XPHY__TXRX_LOOPBACK_5_SZ 40

`define XPHY__TX_DATA_WIDTH    32'h00000047
`define XPHY__TX_DATA_WIDTH_SZ 4

`define XPHY__TX_GATING    32'h00000048
`define XPHY__TX_GATING_SZ 56

`define XPHY__TX_INIT_0    32'h00000049
`define XPHY__TX_INIT_0_SZ 1

`define XPHY__TX_INIT_1    32'h0000004a
`define XPHY__TX_INIT_1_SZ 1

`define XPHY__TX_INIT_2    32'h0000004b
`define XPHY__TX_INIT_2_SZ 1

`define XPHY__TX_INIT_3    32'h0000004c
`define XPHY__TX_INIT_3_SZ 1

`define XPHY__TX_INIT_4    32'h0000004d
`define XPHY__TX_INIT_4_SZ 1

`define XPHY__TX_INIT_5    32'h0000004e
`define XPHY__TX_INIT_5_SZ 1

`define XPHY__TX_INIT_TRI    32'h0000004f
`define XPHY__TX_INIT_TRI_SZ 1

`define XPHY__TX_OUTPUT_PHASE_90_0    32'h00000050
`define XPHY__TX_OUTPUT_PHASE_90_0_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_1    32'h00000051
`define XPHY__TX_OUTPUT_PHASE_90_1_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_2    32'h00000052
`define XPHY__TX_OUTPUT_PHASE_90_2_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_3    32'h00000053
`define XPHY__TX_OUTPUT_PHASE_90_3_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_4    32'h00000054
`define XPHY__TX_OUTPUT_PHASE_90_4_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_5    32'h00000055
`define XPHY__TX_OUTPUT_PHASE_90_5_SZ 40

`define XPHY__TX_OUTPUT_PHASE_90_TRI    32'h00000056
`define XPHY__TX_OUTPUT_PHASE_90_TRI_SZ 40

`define XPHY__WRITE_LEVELING    32'h00000057
`define XPHY__WRITE_LEVELING_SZ 40

`endif  // B_XPHY_DEFINES_VH