// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_MULTIPLIER58_DEFINES_VH
`else
`define B_DSP_MULTIPLIER58_DEFINES_VH

// Look-up table parameters
//

`define DSP_MULTIPLIER58_ADDR_N  5
`define DSP_MULTIPLIER58_ADDR_SZ 32
`define DSP_MULTIPLIER58_DATA_SZ 64

// Attribute addresses
//

`define DSP_MULTIPLIER58__AMULTSEL    32'h00000000
`define DSP_MULTIPLIER58__AMULTSEL_SZ 16

`define DSP_MULTIPLIER58__BMULTSEL    32'h00000001
`define DSP_MULTIPLIER58__BMULTSEL_SZ 16

`define DSP_MULTIPLIER58__DSP_MODE    32'h00000002
`define DSP_MULTIPLIER58__DSP_MODE_SZ 48

`define DSP_MULTIPLIER58__LEGACY    32'h00000003
`define DSP_MULTIPLIER58__LEGACY_SZ 40

`define DSP_MULTIPLIER58__USE_MULT    32'h00000004
`define DSP_MULTIPLIER58__USE_MULT_SZ 64

`endif  // B_DSP_MULTIPLIER58_DEFINES_VH