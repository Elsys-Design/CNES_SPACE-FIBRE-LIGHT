-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description : This module implement the skip insertion word function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
  use phy_plus_lane_lib.all;
  use phy_plus_lane_lib.pkg_phy_plus_lane.all;

entity skip_insertion is
   port (
      RST_N                            : in  std_logic;                       --! global reset
      CLK                              : in  std_logic;                       --! Clock generated by GTY IP

      -- From/to lane_ctrl_word_insert
      NEW_DATA_FROM_LCWI               : in  std_logic;                       --! New data Flag
      DATA_TX_FROM_LCWI                : in  std_logic_vector(31 downto 00);  --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_FROM_LCWI         : in  std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character from DATA-LINK layer
      WAIT_SEND_DATA                   : out std_logic;                       --! Flag to indicates that the lane_ctrl_word_insert send a SKIP control word

      -- To manufacturer IP
      DATA_TX_TO_IP                    : out std_logic_vector(31 downto 00);  --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_TO_IP             : out std_logic_vector(03 downto 00);  --! Flags indicates which byte is a K character

      -- TX signals command from/to lane_init_fsm
      ENABLE_TRANSM_DATA               : in  std_logic                        --! Flag to enable to send data
   );
end skip_insertion;

architecture rtl of skip_insertion is
----------------------------- Declaration signals -----------------------------

signal words_x5000_cnt              : unsigned(12 downto 00);                 --! Allows to count the number of word sent
signal new_data_from_tcwi_r         : std_logic;                              --! NEW_DATA_FROM_LCWI registered signal

begin
-- Send data process
   p_send_data : process(CLK,RST_N)
   begin
      if RST_N = '0' then
         DATA_TX_TO_IP        <= (others => '0');
         VALID_K_CHARAC_TO_IP <= (others => '0');
         words_x5000_cnt      <= (others => '0');
         WAIT_SEND_DATA       <= '0';
         new_data_from_tcwi_r <= '0';

      elsif rising_edge(CLK) then
         new_data_from_tcwi_r <= NEW_DATA_FROM_LCWI;

         if ENABLE_TRANSM_DATA = '1' then                                     -- When the lane_init_fsm is in ACTIVE_ST

            if (NEW_DATA_FROM_LCWI = '1' and new_data_from_tcwi_r = '0') or NEW_DATA_FROM_LCWI = '1' then
               -- Counter 5000 words
               if words_x5000_cnt >= C_5000_WORDS then                        -- When counter reaches 5000
                  WAIT_SEND_DATA       <= '0';                                -- Indicates to the DATA-LINK layer a wait
                  DATA_TX_TO_IP        <= C_SKIP_WORD;                        -- Send SKIP control word
                  VALID_K_CHARAC_TO_IP <= x"1";                               -- Indicates which byte is a K character
                  words_x5000_cnt      <= (others => '0');                    -- Reset counter
               elsif words_x5000_cnt = (C_5000_WORDS -4 )then
                  WAIT_SEND_DATA       <= '1';
                  DATA_TX_TO_IP        <= DATA_TX_FROM_LCWI;                  -- Apply the data fornis by the DATA-LINK layer to the output
                  VALID_K_CHARAC_TO_IP <= VALID_K_CHARAC_FROM_LCWI;           -- Indicates which byte is a K character from DATA-LINK layer
                  words_x5000_cnt      <= words_x5000_cnt+1;  
               elsif words_x5000_cnt < C_5000_WORDS then                      -- else
                  WAIT_SEND_DATA       <= '0';                                -- Indicates the DATA-LINK layer that it can send data
                  DATA_TX_TO_IP        <= DATA_TX_FROM_LCWI;                  -- Apply the data fornis by the DATA-LINK layer to the output
                  VALID_K_CHARAC_TO_IP <= VALID_K_CHARAC_FROM_LCWI;           -- Indicates which byte is a K character from DATA-LINK layer
                  words_x5000_cnt      <= words_x5000_cnt+1;                  -- Increment counter by 1
               end if;
            end if;

         else
            DATA_TX_TO_IP        <= DATA_TX_FROM_LCWI;                        -- Transmit data
            VALID_K_CHARAC_TO_IP <= VALID_K_CHARAC_FROM_LCWI;                 -- Transmit valid K character
            WAIT_SEND_DATA       <= '0';                                      -- And reset all counters and flags
            words_x5000_cnt      <= (others => '0');
         end if;

      end if;
   end process p_send_data;

end architecture rtl;
