`include "B_IOBUFE3_defines.vh"

reg [`IOBUFE3_DATA_SZ-1:0] ATTR [0:`IOBUFE3_ADDR_N-1];
reg [`IOBUFE3__DRIVE_SZ-1:0] DRIVE_REG = DRIVE;
reg [`IOBUFE3__IBUF_LOW_PWR_SZ:1] IBUF_LOW_PWR_REG = IBUF_LOW_PWR;
reg [`IOBUFE3__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IOBUFE3__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`IOBUFE3__SIM_INPUT_BUFFER_OFFSET_SZ-1:0] SIM_INPUT_BUFFER_OFFSET_REG = SIM_INPUT_BUFFER_OFFSET;
reg [`IOBUFE3__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IOBUFE3__DRIVE] = DRIVE;
  ATTR[`IOBUFE3__IBUF_LOW_PWR] = IBUF_LOW_PWR;
  ATTR[`IOBUFE3__IOSTANDARD] = IOSTANDARD;
  ATTR[`IOBUFE3__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`IOBUFE3__SIM_INPUT_BUFFER_OFFSET] = SIM_INPUT_BUFFER_OFFSET;
  ATTR[`IOBUFE3__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  DRIVE_REG = ATTR[`IOBUFE3__DRIVE];
  IBUF_LOW_PWR_REG = ATTR[`IOBUFE3__IBUF_LOW_PWR];
  IOSTANDARD_REG = ATTR[`IOBUFE3__IOSTANDARD];
  SIM_DEVICE_REG = ATTR[`IOBUFE3__SIM_DEVICE];
  SIM_INPUT_BUFFER_OFFSET_REG = ATTR[`IOBUFE3__SIM_INPUT_BUFFER_OFFSET];
  USE_IBUFDISABLE_REG = ATTR[`IOBUFE3__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IOBUFE3_ADDR_SZ-1:0] addr;
  input  [`IOBUFE3_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IOBUFE3_DATA_SZ-1:0] read_attr;
  input  [`IOBUFE3_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
