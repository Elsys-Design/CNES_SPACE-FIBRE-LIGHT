// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_PHY_CHNL_DEFINES_VH
`else
`define B_HBM_PHY_CHNL_DEFINES_VH

// Look-up table parameters
//

`define HBM_PHY_CHNL_ADDR_N  150
`define HBM_PHY_CHNL_ADDR_SZ 32
`define HBM_PHY_CHNL_DATA_SZ 32

// Attribute addresses
//

`define HBM_PHY_CHNL__CFG_00    32'h00000000
`define HBM_PHY_CHNL__CFG_00_SZ 32

`define HBM_PHY_CHNL__CFG_01    32'h00000001
`define HBM_PHY_CHNL__CFG_01_SZ 32

`define HBM_PHY_CHNL__CFG_02    32'h00000002
`define HBM_PHY_CHNL__CFG_02_SZ 31

`define HBM_PHY_CHNL__CFG_03    32'h00000003
`define HBM_PHY_CHNL__CFG_03_SZ 7

`define HBM_PHY_CHNL__CFG_04    32'h00000004
`define HBM_PHY_CHNL__CFG_04_SZ 18

`define HBM_PHY_CHNL__CFG_05    32'h00000005
`define HBM_PHY_CHNL__CFG_05_SZ 18

`define HBM_PHY_CHNL__CFG_06    32'h00000006
`define HBM_PHY_CHNL__CFG_06_SZ 1

`define HBM_PHY_CHNL__CFG_07    32'h00000007
`define HBM_PHY_CHNL__CFG_07_SZ 3

`define HBM_PHY_CHNL__CFG_08    32'h00000008
`define HBM_PHY_CHNL__CFG_08_SZ 32

`define HBM_PHY_CHNL__CFG_09    32'h00000009
`define HBM_PHY_CHNL__CFG_09_SZ 5

`define HBM_PHY_CHNL__CFG_10    32'h0000000a
`define HBM_PHY_CHNL__CFG_10_SZ 11

`define HBM_PHY_CHNL__CFG_100    32'h0000000b
`define HBM_PHY_CHNL__CFG_100_SZ 32

`define HBM_PHY_CHNL__CFG_101    32'h0000000c
`define HBM_PHY_CHNL__CFG_101_SZ 32

`define HBM_PHY_CHNL__CFG_102    32'h0000000d
`define HBM_PHY_CHNL__CFG_102_SZ 32

`define HBM_PHY_CHNL__CFG_103    32'h0000000e
`define HBM_PHY_CHNL__CFG_103_SZ 32

`define HBM_PHY_CHNL__CFG_104    32'h0000000f
`define HBM_PHY_CHNL__CFG_104_SZ 32

`define HBM_PHY_CHNL__CFG_105    32'h00000010
`define HBM_PHY_CHNL__CFG_105_SZ 32

`define HBM_PHY_CHNL__CFG_106    32'h00000011
`define HBM_PHY_CHNL__CFG_106_SZ 32

`define HBM_PHY_CHNL__CFG_107    32'h00000012
`define HBM_PHY_CHNL__CFG_107_SZ 32

`define HBM_PHY_CHNL__CFG_108    32'h00000013
`define HBM_PHY_CHNL__CFG_108_SZ 32

`define HBM_PHY_CHNL__CFG_109    32'h00000014
`define HBM_PHY_CHNL__CFG_109_SZ 32

`define HBM_PHY_CHNL__CFG_11    32'h00000015
`define HBM_PHY_CHNL__CFG_11_SZ 9

`define HBM_PHY_CHNL__CFG_110    32'h00000016
`define HBM_PHY_CHNL__CFG_110_SZ 32

`define HBM_PHY_CHNL__CFG_111    32'h00000017
`define HBM_PHY_CHNL__CFG_111_SZ 9

`define HBM_PHY_CHNL__CFG_112    32'h00000018
`define HBM_PHY_CHNL__CFG_112_SZ 20

`define HBM_PHY_CHNL__CFG_113    32'h00000019
`define HBM_PHY_CHNL__CFG_113_SZ 26

`define HBM_PHY_CHNL__CFG_114    32'h0000001a
`define HBM_PHY_CHNL__CFG_114_SZ 32

`define HBM_PHY_CHNL__CFG_115    32'h0000001b
`define HBM_PHY_CHNL__CFG_115_SZ 6

`define HBM_PHY_CHNL__CFG_116    32'h0000001c
`define HBM_PHY_CHNL__CFG_116_SZ 24

`define HBM_PHY_CHNL__CFG_117    32'h0000001d
`define HBM_PHY_CHNL__CFG_117_SZ 24

`define HBM_PHY_CHNL__CFG_118    32'h0000001e
`define HBM_PHY_CHNL__CFG_118_SZ 24

`define HBM_PHY_CHNL__CFG_119    32'h0000001f
`define HBM_PHY_CHNL__CFG_119_SZ 24

`define HBM_PHY_CHNL__CFG_12    32'h00000020
`define HBM_PHY_CHNL__CFG_12_SZ 13

`define HBM_PHY_CHNL__CFG_120    32'h00000021
`define HBM_PHY_CHNL__CFG_120_SZ 24

`define HBM_PHY_CHNL__CFG_121    32'h00000022
`define HBM_PHY_CHNL__CFG_121_SZ 24

`define HBM_PHY_CHNL__CFG_122    32'h00000023
`define HBM_PHY_CHNL__CFG_122_SZ 24

`define HBM_PHY_CHNL__CFG_123    32'h00000024
`define HBM_PHY_CHNL__CFG_123_SZ 24

`define HBM_PHY_CHNL__CFG_124    32'h00000025
`define HBM_PHY_CHNL__CFG_124_SZ 24

`define HBM_PHY_CHNL__CFG_125    32'h00000026
`define HBM_PHY_CHNL__CFG_125_SZ 24

`define HBM_PHY_CHNL__CFG_126    32'h00000027
`define HBM_PHY_CHNL__CFG_126_SZ 24

`define HBM_PHY_CHNL__CFG_127    32'h00000028
`define HBM_PHY_CHNL__CFG_127_SZ 12

`define HBM_PHY_CHNL__CFG_128    32'h00000029
`define HBM_PHY_CHNL__CFG_128_SZ 12

`define HBM_PHY_CHNL__CFG_129    32'h0000002a
`define HBM_PHY_CHNL__CFG_129_SZ 12

`define HBM_PHY_CHNL__CFG_13    32'h0000002b
`define HBM_PHY_CHNL__CFG_13_SZ 32

`define HBM_PHY_CHNL__CFG_130    32'h0000002c
`define HBM_PHY_CHNL__CFG_130_SZ 23

`define HBM_PHY_CHNL__CFG_131    32'h0000002d
`define HBM_PHY_CHNL__CFG_131_SZ 1

`define HBM_PHY_CHNL__CFG_132    32'h0000002e
`define HBM_PHY_CHNL__CFG_132_SZ 22

`define HBM_PHY_CHNL__CFG_133    32'h0000002f
`define HBM_PHY_CHNL__CFG_133_SZ 23

`define HBM_PHY_CHNL__CFG_134    32'h00000030
`define HBM_PHY_CHNL__CFG_134_SZ 32

`define HBM_PHY_CHNL__CFG_135    32'h00000031
`define HBM_PHY_CHNL__CFG_135_SZ 32

`define HBM_PHY_CHNL__CFG_136    32'h00000032
`define HBM_PHY_CHNL__CFG_136_SZ 32

`define HBM_PHY_CHNL__CFG_137    32'h00000033
`define HBM_PHY_CHNL__CFG_137_SZ 32

`define HBM_PHY_CHNL__CFG_138    32'h00000034
`define HBM_PHY_CHNL__CFG_138_SZ 32

`define HBM_PHY_CHNL__CFG_139    32'h00000035
`define HBM_PHY_CHNL__CFG_139_SZ 32

`define HBM_PHY_CHNL__CFG_14    32'h00000036
`define HBM_PHY_CHNL__CFG_14_SZ 32

`define HBM_PHY_CHNL__CFG_140    32'h00000037
`define HBM_PHY_CHNL__CFG_140_SZ 32

`define HBM_PHY_CHNL__CFG_141    32'h00000038
`define HBM_PHY_CHNL__CFG_141_SZ 32

`define HBM_PHY_CHNL__CFG_142    32'h00000039
`define HBM_PHY_CHNL__CFG_142_SZ 32

`define HBM_PHY_CHNL__CFG_143    32'h0000003a
`define HBM_PHY_CHNL__CFG_143_SZ 24

`define HBM_PHY_CHNL__CFG_144    32'h0000003b
`define HBM_PHY_CHNL__CFG_144_SZ 32

`define HBM_PHY_CHNL__CFG_145    32'h0000003c
`define HBM_PHY_CHNL__CFG_145_SZ 32

`define HBM_PHY_CHNL__CFG_146    32'h0000003d
`define HBM_PHY_CHNL__CFG_146_SZ 32

`define HBM_PHY_CHNL__CFG_147    32'h0000003e
`define HBM_PHY_CHNL__CFG_147_SZ 32

`define HBM_PHY_CHNL__CFG_148    32'h0000003f
`define HBM_PHY_CHNL__CFG_148_SZ 32

`define HBM_PHY_CHNL__CFG_149    32'h00000040
`define HBM_PHY_CHNL__CFG_149_SZ 24

`define HBM_PHY_CHNL__CFG_15    32'h00000041
`define HBM_PHY_CHNL__CFG_15_SZ 8

`define HBM_PHY_CHNL__CFG_16    32'h00000042
`define HBM_PHY_CHNL__CFG_16_SZ 32

`define HBM_PHY_CHNL__CFG_17    32'h00000043
`define HBM_PHY_CHNL__CFG_17_SZ 32

`define HBM_PHY_CHNL__CFG_18    32'h00000044
`define HBM_PHY_CHNL__CFG_18_SZ 32

`define HBM_PHY_CHNL__CFG_19    32'h00000045
`define HBM_PHY_CHNL__CFG_19_SZ 32

`define HBM_PHY_CHNL__CFG_20    32'h00000046
`define HBM_PHY_CHNL__CFG_20_SZ 32

`define HBM_PHY_CHNL__CFG_21    32'h00000047
`define HBM_PHY_CHNL__CFG_21_SZ 30

`define HBM_PHY_CHNL__CFG_23    32'h00000048
`define HBM_PHY_CHNL__CFG_23_SZ 3

`define HBM_PHY_CHNL__CFG_24    32'h00000049
`define HBM_PHY_CHNL__CFG_24_SZ 2

`define HBM_PHY_CHNL__CFG_25    32'h0000004a
`define HBM_PHY_CHNL__CFG_25_SZ 19

`define HBM_PHY_CHNL__CFG_26    32'h0000004b
`define HBM_PHY_CHNL__CFG_26_SZ 17

`define HBM_PHY_CHNL__CFG_27    32'h0000004c
`define HBM_PHY_CHNL__CFG_27_SZ 25

`define HBM_PHY_CHNL__CFG_28    32'h0000004d
`define HBM_PHY_CHNL__CFG_28_SZ 25

`define HBM_PHY_CHNL__CFG_29    32'h0000004e
`define HBM_PHY_CHNL__CFG_29_SZ 25

`define HBM_PHY_CHNL__CFG_30    32'h0000004f
`define HBM_PHY_CHNL__CFG_30_SZ 25

`define HBM_PHY_CHNL__CFG_31    32'h00000050
`define HBM_PHY_CHNL__CFG_31_SZ 25

`define HBM_PHY_CHNL__CFG_32    32'h00000051
`define HBM_PHY_CHNL__CFG_32_SZ 25

`define HBM_PHY_CHNL__CFG_33    32'h00000052
`define HBM_PHY_CHNL__CFG_33_SZ 25

`define HBM_PHY_CHNL__CFG_34    32'h00000053
`define HBM_PHY_CHNL__CFG_34_SZ 25

`define HBM_PHY_CHNL__CFG_35    32'h00000054
`define HBM_PHY_CHNL__CFG_35_SZ 25

`define HBM_PHY_CHNL__CFG_36    32'h00000055
`define HBM_PHY_CHNL__CFG_36_SZ 25

`define HBM_PHY_CHNL__CFG_37    32'h00000056
`define HBM_PHY_CHNL__CFG_37_SZ 25

`define HBM_PHY_CHNL__CFG_38    32'h00000057
`define HBM_PHY_CHNL__CFG_38_SZ 25

`define HBM_PHY_CHNL__CFG_39    32'h00000058
`define HBM_PHY_CHNL__CFG_39_SZ 25

`define HBM_PHY_CHNL__CFG_40    32'h00000059
`define HBM_PHY_CHNL__CFG_40_SZ 25

`define HBM_PHY_CHNL__CFG_41    32'h0000005a
`define HBM_PHY_CHNL__CFG_41_SZ 25

`define HBM_PHY_CHNL__CFG_42    32'h0000005b
`define HBM_PHY_CHNL__CFG_42_SZ 25

`define HBM_PHY_CHNL__CFG_43    32'h0000005c
`define HBM_PHY_CHNL__CFG_43_SZ 25

`define HBM_PHY_CHNL__CFG_44    32'h0000005d
`define HBM_PHY_CHNL__CFG_44_SZ 25

`define HBM_PHY_CHNL__CFG_45    32'h0000005e
`define HBM_PHY_CHNL__CFG_45_SZ 25

`define HBM_PHY_CHNL__CFG_46    32'h0000005f
`define HBM_PHY_CHNL__CFG_46_SZ 25

`define HBM_PHY_CHNL__CFG_47    32'h00000060
`define HBM_PHY_CHNL__CFG_47_SZ 25

`define HBM_PHY_CHNL__CFG_48    32'h00000061
`define HBM_PHY_CHNL__CFG_48_SZ 25

`define HBM_PHY_CHNL__CFG_49    32'h00000062
`define HBM_PHY_CHNL__CFG_49_SZ 25

`define HBM_PHY_CHNL__CFG_50    32'h00000063
`define HBM_PHY_CHNL__CFG_50_SZ 12

`define HBM_PHY_CHNL__CFG_51    32'h00000064
`define HBM_PHY_CHNL__CFG_51_SZ 12

`define HBM_PHY_CHNL__CFG_52    32'h00000065
`define HBM_PHY_CHNL__CFG_52_SZ 12

`define HBM_PHY_CHNL__CFG_53    32'h00000066
`define HBM_PHY_CHNL__CFG_53_SZ 24

`define HBM_PHY_CHNL__CFG_54    32'h00000067
`define HBM_PHY_CHNL__CFG_54_SZ 13

`define HBM_PHY_CHNL__CFG_55    32'h00000068
`define HBM_PHY_CHNL__CFG_55_SZ 10

`define HBM_PHY_CHNL__CFG_56    32'h00000069
`define HBM_PHY_CHNL__CFG_56_SZ 17

`define HBM_PHY_CHNL__CFG_57    32'h0000006a
`define HBM_PHY_CHNL__CFG_57_SZ 8

`define HBM_PHY_CHNL__CFG_58    32'h0000006b
`define HBM_PHY_CHNL__CFG_58_SZ 5

`define HBM_PHY_CHNL__CFG_59    32'h0000006c
`define HBM_PHY_CHNL__CFG_59_SZ 5

`define HBM_PHY_CHNL__CFG_60    32'h0000006d
`define HBM_PHY_CHNL__CFG_60_SZ 16

`define HBM_PHY_CHNL__CFG_61    32'h0000006e
`define HBM_PHY_CHNL__CFG_61_SZ 16

`define HBM_PHY_CHNL__CFG_62    32'h0000006f
`define HBM_PHY_CHNL__CFG_62_SZ 16

`define HBM_PHY_CHNL__CFG_63    32'h00000070
`define HBM_PHY_CHNL__CFG_63_SZ 16

`define HBM_PHY_CHNL__CFG_64    32'h00000071
`define HBM_PHY_CHNL__CFG_64_SZ 20

`define HBM_PHY_CHNL__CFG_65    32'h00000072
`define HBM_PHY_CHNL__CFG_65_SZ 24

`define HBM_PHY_CHNL__CFG_66    32'h00000073
`define HBM_PHY_CHNL__CFG_66_SZ 24

`define HBM_PHY_CHNL__CFG_67    32'h00000074
`define HBM_PHY_CHNL__CFG_67_SZ 32

`define HBM_PHY_CHNL__CFG_68    32'h00000075
`define HBM_PHY_CHNL__CFG_68_SZ 32

`define HBM_PHY_CHNL__CFG_69    32'h00000076
`define HBM_PHY_CHNL__CFG_69_SZ 32

`define HBM_PHY_CHNL__CFG_70    32'h00000077
`define HBM_PHY_CHNL__CFG_70_SZ 32

`define HBM_PHY_CHNL__CFG_71    32'h00000078
`define HBM_PHY_CHNL__CFG_71_SZ 32

`define HBM_PHY_CHNL__CFG_72    32'h00000079
`define HBM_PHY_CHNL__CFG_72_SZ 32

`define HBM_PHY_CHNL__CFG_73    32'h0000007a
`define HBM_PHY_CHNL__CFG_73_SZ 32

`define HBM_PHY_CHNL__CFG_74    32'h0000007b
`define HBM_PHY_CHNL__CFG_74_SZ 32

`define HBM_PHY_CHNL__CFG_75    32'h0000007c
`define HBM_PHY_CHNL__CFG_75_SZ 32

`define HBM_PHY_CHNL__CFG_76    32'h0000007d
`define HBM_PHY_CHNL__CFG_76_SZ 32

`define HBM_PHY_CHNL__CFG_77    32'h0000007e
`define HBM_PHY_CHNL__CFG_77_SZ 32

`define HBM_PHY_CHNL__CFG_78    32'h0000007f
`define HBM_PHY_CHNL__CFG_78_SZ 32

`define HBM_PHY_CHNL__CFG_79    32'h00000080
`define HBM_PHY_CHNL__CFG_79_SZ 32

`define HBM_PHY_CHNL__CFG_80    32'h00000081
`define HBM_PHY_CHNL__CFG_80_SZ 32

`define HBM_PHY_CHNL__CFG_81    32'h00000082
`define HBM_PHY_CHNL__CFG_81_SZ 32

`define HBM_PHY_CHNL__CFG_82    32'h00000083
`define HBM_PHY_CHNL__CFG_82_SZ 32

`define HBM_PHY_CHNL__CFG_83    32'h00000084
`define HBM_PHY_CHNL__CFG_83_SZ 32

`define HBM_PHY_CHNL__CFG_84    32'h00000085
`define HBM_PHY_CHNL__CFG_84_SZ 32

`define HBM_PHY_CHNL__CFG_85    32'h00000086
`define HBM_PHY_CHNL__CFG_85_SZ 16

`define HBM_PHY_CHNL__CFG_86    32'h00000087
`define HBM_PHY_CHNL__CFG_86_SZ 32

`define HBM_PHY_CHNL__CFG_87    32'h00000088
`define HBM_PHY_CHNL__CFG_87_SZ 32

`define HBM_PHY_CHNL__CFG_88    32'h00000089
`define HBM_PHY_CHNL__CFG_88_SZ 4

`define HBM_PHY_CHNL__CFG_89    32'h0000008a
`define HBM_PHY_CHNL__CFG_89_SZ 32

`define HBM_PHY_CHNL__CFG_90    32'h0000008b
`define HBM_PHY_CHNL__CFG_90_SZ 32

`define HBM_PHY_CHNL__CFG_91    32'h0000008c
`define HBM_PHY_CHNL__CFG_91_SZ 24

`define HBM_PHY_CHNL__CFG_92    32'h0000008d
`define HBM_PHY_CHNL__CFG_92_SZ 20

`define HBM_PHY_CHNL__CFG_93    32'h0000008e
`define HBM_PHY_CHNL__CFG_93_SZ 32

`define HBM_PHY_CHNL__CFG_94    32'h0000008f
`define HBM_PHY_CHNL__CFG_94_SZ 32

`define HBM_PHY_CHNL__CFG_95    32'h00000090
`define HBM_PHY_CHNL__CFG_95_SZ 32

`define HBM_PHY_CHNL__CFG_96    32'h00000091
`define HBM_PHY_CHNL__CFG_96_SZ 32

`define HBM_PHY_CHNL__CFG_97    32'h00000092
`define HBM_PHY_CHNL__CFG_97_SZ 32

`define HBM_PHY_CHNL__CFG_98    32'h00000093
`define HBM_PHY_CHNL__CFG_98_SZ 32

`define HBM_PHY_CHNL__CFG_99    32'h00000094
`define HBM_PHY_CHNL__CFG_99_SZ 32

`define HBM_PHY_CHNL__SIM_MODEL_TYPE    32'h00000095
`define HBM_PHY_CHNL__SIM_MODEL_TYPE_SZ 24

`endif  // B_HBM_PHY_CHNL_DEFINES_VH