// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_TX_BITSLICE_TRI_DEFINES_VH
`else
`define B_TX_BITSLICE_TRI_DEFINES_VH

// Look-up table parameters
//

`define TX_BITSLICE_TRI_ADDR_N  14
`define TX_BITSLICE_TRI_ADDR_SZ 32
`define TX_BITSLICE_TRI_DATA_SZ 152

// Attribute addresses
//

`define TX_BITSLICE_TRI__DATA_WIDTH    32'h00000000
`define TX_BITSLICE_TRI__DATA_WIDTH_SZ 4

`define TX_BITSLICE_TRI__DELAY_FORMAT    32'h00000001
`define TX_BITSLICE_TRI__DELAY_FORMAT_SZ 40

`define TX_BITSLICE_TRI__DELAY_TYPE    32'h00000002
`define TX_BITSLICE_TRI__DELAY_TYPE_SZ 64

`define TX_BITSLICE_TRI__DELAY_VALUE    32'h00000003
`define TX_BITSLICE_TRI__DELAY_VALUE_SZ 11

`define TX_BITSLICE_TRI__INIT    32'h00000004
`define TX_BITSLICE_TRI__INIT_SZ 1

`define TX_BITSLICE_TRI__IS_CLK_INVERTED    32'h00000005
`define TX_BITSLICE_TRI__IS_CLK_INVERTED_SZ 1

`define TX_BITSLICE_TRI__IS_RST_DLY_INVERTED    32'h00000006
`define TX_BITSLICE_TRI__IS_RST_DLY_INVERTED_SZ 1

`define TX_BITSLICE_TRI__IS_RST_INVERTED    32'h00000007
`define TX_BITSLICE_TRI__IS_RST_INVERTED_SZ 1

`define TX_BITSLICE_TRI__NATIVE_ODELAY_BYPASS    32'h00000008
`define TX_BITSLICE_TRI__NATIVE_ODELAY_BYPASS_SZ 40

`define TX_BITSLICE_TRI__OUTPUT_PHASE_90    32'h00000009
`define TX_BITSLICE_TRI__OUTPUT_PHASE_90_SZ 40

`define TX_BITSLICE_TRI__REFCLK_FREQUENCY    32'h0000000a
`define TX_BITSLICE_TRI__REFCLK_FREQUENCY_SZ 64

`define TX_BITSLICE_TRI__SIM_DEVICE    32'h0000000b
`define TX_BITSLICE_TRI__SIM_DEVICE_SZ 152

`define TX_BITSLICE_TRI__SIM_VERSION    32'h0000000c
`define TX_BITSLICE_TRI__SIM_VERSION_SZ 64

`define TX_BITSLICE_TRI__UPDATE_MODE    32'h0000000d
`define TX_BITSLICE_TRI__UPDATE_MODE_SZ 48

`endif  // B_TX_BITSLICE_TRI_DEFINES_VH