// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_SYSMONE4_DEFINES_VH
`else
`define B_SYSMONE4_DEFINES_VH

// Look-up table parameters
//

`define SYSMONE4_ADDR_N  77
`define SYSMONE4_ADDR_SZ 32
`define SYSMONE4_DATA_SZ 152

// Attribute addresses
//

`define SYSMONE4__COMMON_N_SOURCE    32'h00000000
`define SYSMONE4__COMMON_N_SOURCE_SZ 16

`define SYSMONE4__INIT_40    32'h00000001
`define SYSMONE4__INIT_40_SZ 16

`define SYSMONE4__INIT_41    32'h00000002
`define SYSMONE4__INIT_41_SZ 16

`define SYSMONE4__INIT_42    32'h00000003
`define SYSMONE4__INIT_42_SZ 16

`define SYSMONE4__INIT_43    32'h00000004
`define SYSMONE4__INIT_43_SZ 16

`define SYSMONE4__INIT_44    32'h00000005
`define SYSMONE4__INIT_44_SZ 16

`define SYSMONE4__INIT_45    32'h00000006
`define SYSMONE4__INIT_45_SZ 16

`define SYSMONE4__INIT_46    32'h00000007
`define SYSMONE4__INIT_46_SZ 16

`define SYSMONE4__INIT_47    32'h00000008
`define SYSMONE4__INIT_47_SZ 16

`define SYSMONE4__INIT_48    32'h00000009
`define SYSMONE4__INIT_48_SZ 16

`define SYSMONE4__INIT_49    32'h0000000a
`define SYSMONE4__INIT_49_SZ 16

`define SYSMONE4__INIT_4A    32'h0000000b
`define SYSMONE4__INIT_4A_SZ 16

`define SYSMONE4__INIT_4B    32'h0000000c
`define SYSMONE4__INIT_4B_SZ 16

`define SYSMONE4__INIT_4C    32'h0000000d
`define SYSMONE4__INIT_4C_SZ 16

`define SYSMONE4__INIT_4D    32'h0000000e
`define SYSMONE4__INIT_4D_SZ 16

`define SYSMONE4__INIT_4E    32'h0000000f
`define SYSMONE4__INIT_4E_SZ 16

`define SYSMONE4__INIT_4F    32'h00000010
`define SYSMONE4__INIT_4F_SZ 16

`define SYSMONE4__INIT_50    32'h00000011
`define SYSMONE4__INIT_50_SZ 16

`define SYSMONE4__INIT_51    32'h00000012
`define SYSMONE4__INIT_51_SZ 16

`define SYSMONE4__INIT_52    32'h00000013
`define SYSMONE4__INIT_52_SZ 16

`define SYSMONE4__INIT_53    32'h00000014
`define SYSMONE4__INIT_53_SZ 16

`define SYSMONE4__INIT_54    32'h00000015
`define SYSMONE4__INIT_54_SZ 16

`define SYSMONE4__INIT_55    32'h00000016
`define SYSMONE4__INIT_55_SZ 16

`define SYSMONE4__INIT_56    32'h00000017
`define SYSMONE4__INIT_56_SZ 16

`define SYSMONE4__INIT_57    32'h00000018
`define SYSMONE4__INIT_57_SZ 16

`define SYSMONE4__INIT_58    32'h00000019
`define SYSMONE4__INIT_58_SZ 16

`define SYSMONE4__INIT_59    32'h0000001a
`define SYSMONE4__INIT_59_SZ 16

`define SYSMONE4__INIT_5A    32'h0000001b
`define SYSMONE4__INIT_5A_SZ 16

`define SYSMONE4__INIT_5B    32'h0000001c
`define SYSMONE4__INIT_5B_SZ 16

`define SYSMONE4__INIT_5C    32'h0000001d
`define SYSMONE4__INIT_5C_SZ 16

`define SYSMONE4__INIT_5D    32'h0000001e
`define SYSMONE4__INIT_5D_SZ 16

`define SYSMONE4__INIT_5E    32'h0000001f
`define SYSMONE4__INIT_5E_SZ 16

`define SYSMONE4__INIT_5F    32'h00000020
`define SYSMONE4__INIT_5F_SZ 16

`define SYSMONE4__INIT_60    32'h00000021
`define SYSMONE4__INIT_60_SZ 16

`define SYSMONE4__INIT_61    32'h00000022
`define SYSMONE4__INIT_61_SZ 16

`define SYSMONE4__INIT_62    32'h00000023
`define SYSMONE4__INIT_62_SZ 16

`define SYSMONE4__INIT_63    32'h00000024
`define SYSMONE4__INIT_63_SZ 16

`define SYSMONE4__INIT_64    32'h00000025
`define SYSMONE4__INIT_64_SZ 16

`define SYSMONE4__INIT_65    32'h00000026
`define SYSMONE4__INIT_65_SZ 16

`define SYSMONE4__INIT_66    32'h00000027
`define SYSMONE4__INIT_66_SZ 16

`define SYSMONE4__INIT_67    32'h00000028
`define SYSMONE4__INIT_67_SZ 16

`define SYSMONE4__INIT_68    32'h00000029
`define SYSMONE4__INIT_68_SZ 16

`define SYSMONE4__INIT_69    32'h0000002a
`define SYSMONE4__INIT_69_SZ 16

`define SYSMONE4__INIT_6A    32'h0000002b
`define SYSMONE4__INIT_6A_SZ 16

`define SYSMONE4__INIT_6B    32'h0000002c
`define SYSMONE4__INIT_6B_SZ 16

`define SYSMONE4__INIT_6C    32'h0000002d
`define SYSMONE4__INIT_6C_SZ 16

`define SYSMONE4__INIT_6D    32'h0000002e
`define SYSMONE4__INIT_6D_SZ 16

`define SYSMONE4__INIT_6E    32'h0000002f
`define SYSMONE4__INIT_6E_SZ 16

`define SYSMONE4__INIT_6F    32'h00000030
`define SYSMONE4__INIT_6F_SZ 16

`define SYSMONE4__INIT_70    32'h00000031
`define SYSMONE4__INIT_70_SZ 16

`define SYSMONE4__INIT_71    32'h00000032
`define SYSMONE4__INIT_71_SZ 16

`define SYSMONE4__INIT_72    32'h00000033
`define SYSMONE4__INIT_72_SZ 16

`define SYSMONE4__INIT_73    32'h00000034
`define SYSMONE4__INIT_73_SZ 16

`define SYSMONE4__INIT_74    32'h00000035
`define SYSMONE4__INIT_74_SZ 16

`define SYSMONE4__INIT_75    32'h00000036
`define SYSMONE4__INIT_75_SZ 16

`define SYSMONE4__INIT_76    32'h00000037
`define SYSMONE4__INIT_76_SZ 16

`define SYSMONE4__INIT_77    32'h00000038
`define SYSMONE4__INIT_77_SZ 16

`define SYSMONE4__INIT_78    32'h00000039
`define SYSMONE4__INIT_78_SZ 16

`define SYSMONE4__INIT_79    32'h0000003a
`define SYSMONE4__INIT_79_SZ 16

`define SYSMONE4__INIT_7A    32'h0000003b
`define SYSMONE4__INIT_7A_SZ 16

`define SYSMONE4__INIT_7B    32'h0000003c
`define SYSMONE4__INIT_7B_SZ 16

`define SYSMONE4__INIT_7C    32'h0000003d
`define SYSMONE4__INIT_7C_SZ 16

`define SYSMONE4__INIT_7D    32'h0000003e
`define SYSMONE4__INIT_7D_SZ 16

`define SYSMONE4__INIT_7E    32'h0000003f
`define SYSMONE4__INIT_7E_SZ 16

`define SYSMONE4__INIT_7F    32'h00000040
`define SYSMONE4__INIT_7F_SZ 16

`define SYSMONE4__IS_CONVSTCLK_INVERTED    32'h00000041
`define SYSMONE4__IS_CONVSTCLK_INVERTED_SZ 1

`define SYSMONE4__IS_DCLK_INVERTED    32'h00000042
`define SYSMONE4__IS_DCLK_INVERTED_SZ 1

`define SYSMONE4__SIM_DEVICE    32'h00000043
`define SYSMONE4__SIM_DEVICE_SZ 152

`define SYSMONE4__SIM_MONITOR_FILE    32'h00000044
`define SYSMONE4__SIM_MONITOR_FILE_SZ 80

`define SYSMONE4__SYSMON_VUSER0_BANK    32'h00000045
`define SYSMONE4__SYSMON_VUSER0_BANK_SZ 32

`define SYSMONE4__SYSMON_VUSER0_MONITOR    32'h00000046
`define SYSMONE4__SYSMON_VUSER0_MONITOR_SZ 32

`define SYSMONE4__SYSMON_VUSER1_BANK    32'h00000047
`define SYSMONE4__SYSMON_VUSER1_BANK_SZ 32

`define SYSMONE4__SYSMON_VUSER1_MONITOR    32'h00000048
`define SYSMONE4__SYSMON_VUSER1_MONITOR_SZ 32

`define SYSMONE4__SYSMON_VUSER2_BANK    32'h00000049
`define SYSMONE4__SYSMON_VUSER2_BANK_SZ 32

`define SYSMONE4__SYSMON_VUSER2_MONITOR    32'h0000004a
`define SYSMONE4__SYSMON_VUSER2_MONITOR_SZ 32

`define SYSMONE4__SYSMON_VUSER3_BANK    32'h0000004b
`define SYSMONE4__SYSMON_VUSER3_BANK_SZ 32

`define SYSMONE4__SYSMON_VUSER3_MONITOR    32'h0000004c
`define SYSMONE4__SYSMON_VUSER3_MONITOR_SZ 32

`endif  // B_SYSMONE4_DEFINES_VH