// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_MRMAC_DEFINES_VH
`else
`define B_MRMAC_DEFINES_VH

// Look-up table parameters
//

`define MRMAC_ADDR_N  568
`define MRMAC_ADDR_SZ 32
`define MRMAC_DATA_SZ 144

// Attribute addresses
//

`define MRMAC__ACTIVITY    32'h00000000
`define MRMAC__ACTIVITY_SZ 56

`define MRMAC__CTL_AXIS_CFG_0    32'h00000001
`define MRMAC__CTL_AXIS_CFG_0_SZ 3

`define MRMAC__CTL_AXIS_CFG_1    32'h00000002
`define MRMAC__CTL_AXIS_CFG_1_SZ 3

`define MRMAC__CTL_AXIS_CFG_2    32'h00000003
`define MRMAC__CTL_AXIS_CFG_2_SZ 3

`define MRMAC__CTL_AXIS_CFG_3    32'h00000004
`define MRMAC__CTL_AXIS_CFG_3_SZ 3

`define MRMAC__CTL_COUNTER_EXTEND_0    32'h00000005
`define MRMAC__CTL_COUNTER_EXTEND_0_SZ 40

`define MRMAC__CTL_COUNTER_EXTEND_1    32'h00000006
`define MRMAC__CTL_COUNTER_EXTEND_1_SZ 40

`define MRMAC__CTL_COUNTER_EXTEND_2    32'h00000007
`define MRMAC__CTL_COUNTER_EXTEND_2_SZ 40

`define MRMAC__CTL_COUNTER_EXTEND_3    32'h00000008
`define MRMAC__CTL_COUNTER_EXTEND_3_SZ 40

`define MRMAC__CTL_CUSTOM_RX_AMS_0    32'h00000009
`define MRMAC__CTL_CUSTOM_RX_AMS_0_SZ 40

`define MRMAC__CTL_CUSTOM_RX_AMS_1    32'h0000000a
`define MRMAC__CTL_CUSTOM_RX_AMS_1_SZ 40

`define MRMAC__CTL_CUSTOM_RX_AMS_2    32'h0000000b
`define MRMAC__CTL_CUSTOM_RX_AMS_2_SZ 40

`define MRMAC__CTL_CUSTOM_RX_AMS_3    32'h0000000c
`define MRMAC__CTL_CUSTOM_RX_AMS_3_SZ 40

`define MRMAC__CTL_CUSTOM_TX_AMS_0    32'h0000000d
`define MRMAC__CTL_CUSTOM_TX_AMS_0_SZ 40

`define MRMAC__CTL_CUSTOM_TX_AMS_1    32'h0000000e
`define MRMAC__CTL_CUSTOM_TX_AMS_1_SZ 40

`define MRMAC__CTL_CUSTOM_TX_AMS_2    32'h0000000f
`define MRMAC__CTL_CUSTOM_TX_AMS_2_SZ 40

`define MRMAC__CTL_CUSTOM_TX_AMS_3    32'h00000010
`define MRMAC__CTL_CUSTOM_TX_AMS_3_SZ 40

`define MRMAC__CTL_DATA_RATE_0    32'h00000011
`define MRMAC__CTL_DATA_RATE_0_SZ 3

`define MRMAC__CTL_DATA_RATE_1    32'h00000012
`define MRMAC__CTL_DATA_RATE_1_SZ 2

`define MRMAC__CTL_DATA_RATE_2    32'h00000013
`define MRMAC__CTL_DATA_RATE_2_SZ 2

`define MRMAC__CTL_DATA_RATE_3    32'h00000014
`define MRMAC__CTL_DATA_RATE_3_SZ 2

`define MRMAC__CTL_FEC_MODE_0    32'h00000015
`define MRMAC__CTL_FEC_MODE_0_SZ 4

`define MRMAC__CTL_FEC_MODE_1    32'h00000016
`define MRMAC__CTL_FEC_MODE_1_SZ 4

`define MRMAC__CTL_FEC_MODE_2    32'h00000017
`define MRMAC__CTL_FEC_MODE_2_SZ 4

`define MRMAC__CTL_FEC_MODE_3    32'h00000018
`define MRMAC__CTL_FEC_MODE_3_SZ 4

`define MRMAC__CTL_PCS_RX_TS_EN_0    32'h00000019
`define MRMAC__CTL_PCS_RX_TS_EN_0_SZ 40

`define MRMAC__CTL_PCS_RX_TS_EN_1    32'h0000001a
`define MRMAC__CTL_PCS_RX_TS_EN_1_SZ 40

`define MRMAC__CTL_PCS_RX_TS_EN_2    32'h0000001b
`define MRMAC__CTL_PCS_RX_TS_EN_2_SZ 40

`define MRMAC__CTL_PCS_RX_TS_EN_3    32'h0000001c
`define MRMAC__CTL_PCS_RX_TS_EN_3_SZ 40

`define MRMAC__CTL_PREEMPT_ENABLE_0    32'h0000001d
`define MRMAC__CTL_PREEMPT_ENABLE_0_SZ 40

`define MRMAC__CTL_PREEMPT_ENABLE_1    32'h0000001e
`define MRMAC__CTL_PREEMPT_ENABLE_1_SZ 40

`define MRMAC__CTL_PREEMPT_ENABLE_2    32'h0000001f
`define MRMAC__CTL_PREEMPT_ENABLE_2_SZ 40

`define MRMAC__CTL_PREEMPT_ENABLE_3    32'h00000020
`define MRMAC__CTL_PREEMPT_ENABLE_3_SZ 40

`define MRMAC__CTL_REVISION    32'h00000021
`define MRMAC__CTL_REVISION_SZ 32

`define MRMAC__CTL_RX01_DEGRADE_ACT_THRESH    32'h00000022
`define MRMAC__CTL_RX01_DEGRADE_ACT_THRESH_SZ 16

`define MRMAC__CTL_RX01_DEGRADE_DEACT_THRESH    32'h00000023
`define MRMAC__CTL_RX01_DEGRADE_DEACT_THRESH_SZ 16

`define MRMAC__CTL_RX01_DEGRADE_ENABLE    32'h00000024
`define MRMAC__CTL_RX01_DEGRADE_ENABLE_SZ 40

`define MRMAC__CTL_RX01_DEGRADE_INTERVAL    32'h00000025
`define MRMAC__CTL_RX01_DEGRADE_INTERVAL_SZ 16

`define MRMAC__CTL_RX23_DEGRADE_ACT_THRESH    32'h00000026
`define MRMAC__CTL_RX23_DEGRADE_ACT_THRESH_SZ 16

`define MRMAC__CTL_RX23_DEGRADE_DEACT_THRESH    32'h00000027
`define MRMAC__CTL_RX23_DEGRADE_DEACT_THRESH_SZ 16

`define MRMAC__CTL_RX23_DEGRADE_ENABLE    32'h00000028
`define MRMAC__CTL_RX23_DEGRADE_ENABLE_SZ 40

`define MRMAC__CTL_RX23_DEGRADE_INTERVAL    32'h00000029
`define MRMAC__CTL_RX23_DEGRADE_INTERVAL_SZ 16

`define MRMAC__CTL_RX_CHECK_ACK_0    32'h0000002a
`define MRMAC__CTL_RX_CHECK_ACK_0_SZ 40

`define MRMAC__CTL_RX_CHECK_ACK_1    32'h0000002b
`define MRMAC__CTL_RX_CHECK_ACK_1_SZ 40

`define MRMAC__CTL_RX_CHECK_ACK_2    32'h0000002c
`define MRMAC__CTL_RX_CHECK_ACK_2_SZ 40

`define MRMAC__CTL_RX_CHECK_ACK_3    32'h0000002d
`define MRMAC__CTL_RX_CHECK_ACK_3_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_0    32'h0000002e
`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_1    32'h0000002f
`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_2    32'h00000030
`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_3    32'h00000031
`define MRMAC__CTL_RX_CHECK_ETYPE_GCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_0    32'h00000032
`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_1    32'h00000033
`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_2    32'h00000034
`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_3    32'h00000035
`define MRMAC__CTL_RX_CHECK_ETYPE_GPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_0    32'h00000036
`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_1    32'h00000037
`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_2    32'h00000038
`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_3    32'h00000039
`define MRMAC__CTL_RX_CHECK_ETYPE_PCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_0    32'h0000003a
`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_1    32'h0000003b
`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_2    32'h0000003c
`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_3    32'h0000003d
`define MRMAC__CTL_RX_CHECK_ETYPE_PPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GCP_0    32'h0000003e
`define MRMAC__CTL_RX_CHECK_MCAST_GCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GCP_1    32'h0000003f
`define MRMAC__CTL_RX_CHECK_MCAST_GCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GCP_2    32'h00000040
`define MRMAC__CTL_RX_CHECK_MCAST_GCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GCP_3    32'h00000041
`define MRMAC__CTL_RX_CHECK_MCAST_GCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GPP_0    32'h00000042
`define MRMAC__CTL_RX_CHECK_MCAST_GPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GPP_1    32'h00000043
`define MRMAC__CTL_RX_CHECK_MCAST_GPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GPP_2    32'h00000044
`define MRMAC__CTL_RX_CHECK_MCAST_GPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_GPP_3    32'h00000045
`define MRMAC__CTL_RX_CHECK_MCAST_GPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PCP_0    32'h00000046
`define MRMAC__CTL_RX_CHECK_MCAST_PCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PCP_1    32'h00000047
`define MRMAC__CTL_RX_CHECK_MCAST_PCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PCP_2    32'h00000048
`define MRMAC__CTL_RX_CHECK_MCAST_PCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PCP_3    32'h00000049
`define MRMAC__CTL_RX_CHECK_MCAST_PCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PPP_0    32'h0000004a
`define MRMAC__CTL_RX_CHECK_MCAST_PPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PPP_1    32'h0000004b
`define MRMAC__CTL_RX_CHECK_MCAST_PPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PPP_2    32'h0000004c
`define MRMAC__CTL_RX_CHECK_MCAST_PPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_MCAST_PPP_3    32'h0000004d
`define MRMAC__CTL_RX_CHECK_MCAST_PPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_0    32'h0000004e
`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_1    32'h0000004f
`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_2    32'h00000050
`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_3    32'h00000051
`define MRMAC__CTL_RX_CHECK_OPCODE_GCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_0    32'h00000052
`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_1    32'h00000053
`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_2    32'h00000054
`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_3    32'h00000055
`define MRMAC__CTL_RX_CHECK_OPCODE_GPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_0    32'h00000056
`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_1    32'h00000057
`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_2    32'h00000058
`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_3    32'h00000059
`define MRMAC__CTL_RX_CHECK_OPCODE_PCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_0    32'h0000005a
`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_1    32'h0000005b
`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_2    32'h0000005c
`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_3    32'h0000005d
`define MRMAC__CTL_RX_CHECK_OPCODE_PPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_PREAMBLE_0    32'h0000005e
`define MRMAC__CTL_RX_CHECK_PREAMBLE_0_SZ 40

`define MRMAC__CTL_RX_CHECK_PREAMBLE_1    32'h0000005f
`define MRMAC__CTL_RX_CHECK_PREAMBLE_1_SZ 40

`define MRMAC__CTL_RX_CHECK_PREAMBLE_2    32'h00000060
`define MRMAC__CTL_RX_CHECK_PREAMBLE_2_SZ 40

`define MRMAC__CTL_RX_CHECK_PREAMBLE_3    32'h00000061
`define MRMAC__CTL_RX_CHECK_PREAMBLE_3_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GCP_0    32'h00000062
`define MRMAC__CTL_RX_CHECK_SA_GCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GCP_1    32'h00000063
`define MRMAC__CTL_RX_CHECK_SA_GCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GCP_2    32'h00000064
`define MRMAC__CTL_RX_CHECK_SA_GCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GCP_3    32'h00000065
`define MRMAC__CTL_RX_CHECK_SA_GCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GPP_0    32'h00000066
`define MRMAC__CTL_RX_CHECK_SA_GPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GPP_1    32'h00000067
`define MRMAC__CTL_RX_CHECK_SA_GPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GPP_2    32'h00000068
`define MRMAC__CTL_RX_CHECK_SA_GPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_GPP_3    32'h00000069
`define MRMAC__CTL_RX_CHECK_SA_GPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PCP_0    32'h0000006a
`define MRMAC__CTL_RX_CHECK_SA_PCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PCP_1    32'h0000006b
`define MRMAC__CTL_RX_CHECK_SA_PCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PCP_2    32'h0000006c
`define MRMAC__CTL_RX_CHECK_SA_PCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PCP_3    32'h0000006d
`define MRMAC__CTL_RX_CHECK_SA_PCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PPP_0    32'h0000006e
`define MRMAC__CTL_RX_CHECK_SA_PPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PPP_1    32'h0000006f
`define MRMAC__CTL_RX_CHECK_SA_PPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PPP_2    32'h00000070
`define MRMAC__CTL_RX_CHECK_SA_PPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_SA_PPP_3    32'h00000071
`define MRMAC__CTL_RX_CHECK_SA_PPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_SFD_0    32'h00000072
`define MRMAC__CTL_RX_CHECK_SFD_0_SZ 40

`define MRMAC__CTL_RX_CHECK_SFD_1    32'h00000073
`define MRMAC__CTL_RX_CHECK_SFD_1_SZ 40

`define MRMAC__CTL_RX_CHECK_SFD_2    32'h00000074
`define MRMAC__CTL_RX_CHECK_SFD_2_SZ 40

`define MRMAC__CTL_RX_CHECK_SFD_3    32'h00000075
`define MRMAC__CTL_RX_CHECK_SFD_3_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GCP_0    32'h00000076
`define MRMAC__CTL_RX_CHECK_UCAST_GCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GCP_1    32'h00000077
`define MRMAC__CTL_RX_CHECK_UCAST_GCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GCP_2    32'h00000078
`define MRMAC__CTL_RX_CHECK_UCAST_GCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GCP_3    32'h00000079
`define MRMAC__CTL_RX_CHECK_UCAST_GCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GPP_0    32'h0000007a
`define MRMAC__CTL_RX_CHECK_UCAST_GPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GPP_1    32'h0000007b
`define MRMAC__CTL_RX_CHECK_UCAST_GPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GPP_2    32'h0000007c
`define MRMAC__CTL_RX_CHECK_UCAST_GPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_GPP_3    32'h0000007d
`define MRMAC__CTL_RX_CHECK_UCAST_GPP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PCP_0    32'h0000007e
`define MRMAC__CTL_RX_CHECK_UCAST_PCP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PCP_1    32'h0000007f
`define MRMAC__CTL_RX_CHECK_UCAST_PCP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PCP_2    32'h00000080
`define MRMAC__CTL_RX_CHECK_UCAST_PCP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PCP_3    32'h00000081
`define MRMAC__CTL_RX_CHECK_UCAST_PCP_3_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PPP_0    32'h00000082
`define MRMAC__CTL_RX_CHECK_UCAST_PPP_0_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PPP_1    32'h00000083
`define MRMAC__CTL_RX_CHECK_UCAST_PPP_1_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PPP_2    32'h00000084
`define MRMAC__CTL_RX_CHECK_UCAST_PPP_2_SZ 40

`define MRMAC__CTL_RX_CHECK_UCAST_PPP_3    32'h00000085
`define MRMAC__CTL_RX_CHECK_UCAST_PPP_3_SZ 40

`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_0    32'h00000086
`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_0_SZ 40

`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_1    32'h00000087
`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_1_SZ 40

`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_2    32'h00000088
`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_2_SZ 40

`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_3    32'h00000089
`define MRMAC__CTL_RX_DATA_PATTERN_SELECT_3_SZ 40

`define MRMAC__CTL_RX_DELETE_FCS_0    32'h0000008a
`define MRMAC__CTL_RX_DELETE_FCS_0_SZ 40

`define MRMAC__CTL_RX_DELETE_FCS_1    32'h0000008b
`define MRMAC__CTL_RX_DELETE_FCS_1_SZ 40

`define MRMAC__CTL_RX_DELETE_FCS_2    32'h0000008c
`define MRMAC__CTL_RX_DELETE_FCS_2_SZ 40

`define MRMAC__CTL_RX_DELETE_FCS_3    32'h0000008d
`define MRMAC__CTL_RX_DELETE_FCS_3_SZ 40

`define MRMAC__CTL_RX_ENABLE_0    32'h0000008e
`define MRMAC__CTL_RX_ENABLE_0_SZ 40

`define MRMAC__CTL_RX_ENABLE_1    32'h0000008f
`define MRMAC__CTL_RX_ENABLE_1_SZ 40

`define MRMAC__CTL_RX_ENABLE_2    32'h00000090
`define MRMAC__CTL_RX_ENABLE_2_SZ 40

`define MRMAC__CTL_RX_ENABLE_3    32'h00000091
`define MRMAC__CTL_RX_ENABLE_3_SZ 40

`define MRMAC__CTL_RX_ENABLE_GCP_0    32'h00000092
`define MRMAC__CTL_RX_ENABLE_GCP_0_SZ 40

`define MRMAC__CTL_RX_ENABLE_GCP_1    32'h00000093
`define MRMAC__CTL_RX_ENABLE_GCP_1_SZ 40

`define MRMAC__CTL_RX_ENABLE_GCP_2    32'h00000094
`define MRMAC__CTL_RX_ENABLE_GCP_2_SZ 40

`define MRMAC__CTL_RX_ENABLE_GCP_3    32'h00000095
`define MRMAC__CTL_RX_ENABLE_GCP_3_SZ 40

`define MRMAC__CTL_RX_ENABLE_GPP_0    32'h00000096
`define MRMAC__CTL_RX_ENABLE_GPP_0_SZ 40

`define MRMAC__CTL_RX_ENABLE_GPP_1    32'h00000097
`define MRMAC__CTL_RX_ENABLE_GPP_1_SZ 40

`define MRMAC__CTL_RX_ENABLE_GPP_2    32'h00000098
`define MRMAC__CTL_RX_ENABLE_GPP_2_SZ 40

`define MRMAC__CTL_RX_ENABLE_GPP_3    32'h00000099
`define MRMAC__CTL_RX_ENABLE_GPP_3_SZ 40

`define MRMAC__CTL_RX_ENABLE_PCP_0    32'h0000009a
`define MRMAC__CTL_RX_ENABLE_PCP_0_SZ 40

`define MRMAC__CTL_RX_ENABLE_PCP_1    32'h0000009b
`define MRMAC__CTL_RX_ENABLE_PCP_1_SZ 40

`define MRMAC__CTL_RX_ENABLE_PCP_2    32'h0000009c
`define MRMAC__CTL_RX_ENABLE_PCP_2_SZ 40

`define MRMAC__CTL_RX_ENABLE_PCP_3    32'h0000009d
`define MRMAC__CTL_RX_ENABLE_PCP_3_SZ 40

`define MRMAC__CTL_RX_ENABLE_PPP_0    32'h0000009e
`define MRMAC__CTL_RX_ENABLE_PPP_0_SZ 40

`define MRMAC__CTL_RX_ENABLE_PPP_1    32'h0000009f
`define MRMAC__CTL_RX_ENABLE_PPP_1_SZ 40

`define MRMAC__CTL_RX_ENABLE_PPP_2    32'h000000a0
`define MRMAC__CTL_RX_ENABLE_PPP_2_SZ 40

`define MRMAC__CTL_RX_ENABLE_PPP_3    32'h000000a1
`define MRMAC__CTL_RX_ENABLE_PPP_3_SZ 40

`define MRMAC__CTL_RX_ETYPE_GCP_0    32'h000000a2
`define MRMAC__CTL_RX_ETYPE_GCP_0_SZ 16

`define MRMAC__CTL_RX_ETYPE_GCP_1    32'h000000a3
`define MRMAC__CTL_RX_ETYPE_GCP_1_SZ 16

`define MRMAC__CTL_RX_ETYPE_GCP_2    32'h000000a4
`define MRMAC__CTL_RX_ETYPE_GCP_2_SZ 16

`define MRMAC__CTL_RX_ETYPE_GCP_3    32'h000000a5
`define MRMAC__CTL_RX_ETYPE_GCP_3_SZ 16

`define MRMAC__CTL_RX_ETYPE_GPP_0    32'h000000a6
`define MRMAC__CTL_RX_ETYPE_GPP_0_SZ 16

`define MRMAC__CTL_RX_ETYPE_GPP_1    32'h000000a7
`define MRMAC__CTL_RX_ETYPE_GPP_1_SZ 16

`define MRMAC__CTL_RX_ETYPE_GPP_2    32'h000000a8
`define MRMAC__CTL_RX_ETYPE_GPP_2_SZ 16

`define MRMAC__CTL_RX_ETYPE_GPP_3    32'h000000a9
`define MRMAC__CTL_RX_ETYPE_GPP_3_SZ 16

`define MRMAC__CTL_RX_ETYPE_PCP_0    32'h000000aa
`define MRMAC__CTL_RX_ETYPE_PCP_0_SZ 16

`define MRMAC__CTL_RX_ETYPE_PCP_1    32'h000000ab
`define MRMAC__CTL_RX_ETYPE_PCP_1_SZ 16

`define MRMAC__CTL_RX_ETYPE_PCP_2    32'h000000ac
`define MRMAC__CTL_RX_ETYPE_PCP_2_SZ 16

`define MRMAC__CTL_RX_ETYPE_PCP_3    32'h000000ad
`define MRMAC__CTL_RX_ETYPE_PCP_3_SZ 16

`define MRMAC__CTL_RX_ETYPE_PPP_0    32'h000000ae
`define MRMAC__CTL_RX_ETYPE_PPP_0_SZ 16

`define MRMAC__CTL_RX_ETYPE_PPP_1    32'h000000af
`define MRMAC__CTL_RX_ETYPE_PPP_1_SZ 16

`define MRMAC__CTL_RX_ETYPE_PPP_2    32'h000000b0
`define MRMAC__CTL_RX_ETYPE_PPP_2_SZ 16

`define MRMAC__CTL_RX_ETYPE_PPP_3    32'h000000b1
`define MRMAC__CTL_RX_ETYPE_PPP_3_SZ 16

`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_0    32'h000000b2
`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_0_SZ 40

`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_1    32'h000000b3
`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_1_SZ 40

`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_2    32'h000000b4
`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_2_SZ 40

`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_3    32'h000000b5
`define MRMAC__CTL_RX_FEC_ALIGNMENT_BYPASS_3_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_0    32'h000000b6
`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_0_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_1    32'h000000b7
`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_1_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_2    32'h000000b8
`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_2_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_3    32'h000000b9
`define MRMAC__CTL_RX_FEC_BYPASS_CORRECTION_3_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_0    32'h000000ba
`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_0_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_1    32'h000000bb
`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_1_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_2    32'h000000bc
`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_2_SZ 40

`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_3    32'h000000bd
`define MRMAC__CTL_RX_FEC_BYPASS_INDICATION_3_SZ 40

`define MRMAC__CTL_RX_FEC_CDC_BYPASS_01    32'h000000be
`define MRMAC__CTL_RX_FEC_CDC_BYPASS_01_SZ 40

`define MRMAC__CTL_RX_FEC_CDC_BYPASS_23    32'h000000bf
`define MRMAC__CTL_RX_FEC_CDC_BYPASS_23_SZ 40

`define MRMAC__CTL_RX_FEC_ERRIND_MODE    32'h000000c0
`define MRMAC__CTL_RX_FEC_ERRIND_MODE_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_0    32'h000000c1
`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_0_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_1    32'h000000c2
`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_1_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_2    32'h000000c3
`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_2_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_3    32'h000000c4
`define MRMAC__CTL_RX_FEC_TRANSCODE_BYPASS_3_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_0    32'h000000c5
`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_0_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_1    32'h000000c6
`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_1_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_2    32'h000000c7
`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_2_SZ 40

`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_3    32'h000000c8
`define MRMAC__CTL_RX_FEC_TRANSCODE_CLAUSE49_3_SZ 40

`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_0    32'h000000c9
`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_0_SZ 40

`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_1    32'h000000ca
`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_1_SZ 40

`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_2    32'h000000cb
`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_2_SZ 40

`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_3    32'h000000cc
`define MRMAC__CTL_RX_FLEXIF_INPUT_ENABLE_3_SZ 40

`define MRMAC__CTL_RX_FLEXIF_SELECT_0    32'h000000cd
`define MRMAC__CTL_RX_FLEXIF_SELECT_0_SZ 4

`define MRMAC__CTL_RX_FLEXIF_SELECT_1    32'h000000ce
`define MRMAC__CTL_RX_FLEXIF_SELECT_1_SZ 4

`define MRMAC__CTL_RX_FLEXIF_SELECT_2    32'h000000cf
`define MRMAC__CTL_RX_FLEXIF_SELECT_2_SZ 4

`define MRMAC__CTL_RX_FLEXIF_SELECT_3    32'h000000d0
`define MRMAC__CTL_RX_FLEXIF_SELECT_3_SZ 4

`define MRMAC__CTL_RX_FORWARD_CONTROL_0    32'h000000d1
`define MRMAC__CTL_RX_FORWARD_CONTROL_0_SZ 40

`define MRMAC__CTL_RX_FORWARD_CONTROL_1    32'h000000d2
`define MRMAC__CTL_RX_FORWARD_CONTROL_1_SZ 40

`define MRMAC__CTL_RX_FORWARD_CONTROL_2    32'h000000d3
`define MRMAC__CTL_RX_FORWARD_CONTROL_2_SZ 40

`define MRMAC__CTL_RX_FORWARD_CONTROL_3    32'h000000d4
`define MRMAC__CTL_RX_FORWARD_CONTROL_3_SZ 40

`define MRMAC__CTL_RX_IGNORE_FCS_0    32'h000000d5
`define MRMAC__CTL_RX_IGNORE_FCS_0_SZ 40

`define MRMAC__CTL_RX_IGNORE_FCS_1    32'h000000d6
`define MRMAC__CTL_RX_IGNORE_FCS_1_SZ 40

`define MRMAC__CTL_RX_IGNORE_FCS_2    32'h000000d7
`define MRMAC__CTL_RX_IGNORE_FCS_2_SZ 40

`define MRMAC__CTL_RX_IGNORE_FCS_3    32'h000000d8
`define MRMAC__CTL_RX_IGNORE_FCS_3_SZ 40

`define MRMAC__CTL_RX_IGNORE_INRANGE_0    32'h000000d9
`define MRMAC__CTL_RX_IGNORE_INRANGE_0_SZ 40

`define MRMAC__CTL_RX_IGNORE_INRANGE_1    32'h000000da
`define MRMAC__CTL_RX_IGNORE_INRANGE_1_SZ 40

`define MRMAC__CTL_RX_IGNORE_INRANGE_2    32'h000000db
`define MRMAC__CTL_RX_IGNORE_INRANGE_2_SZ 40

`define MRMAC__CTL_RX_IGNORE_INRANGE_3    32'h000000dc
`define MRMAC__CTL_RX_IGNORE_INRANGE_3_SZ 40

`define MRMAC__CTL_RX_MAX_PACKET_LEN_0    32'h000000dd
`define MRMAC__CTL_RX_MAX_PACKET_LEN_0_SZ 15

`define MRMAC__CTL_RX_MAX_PACKET_LEN_1    32'h000000de
`define MRMAC__CTL_RX_MAX_PACKET_LEN_1_SZ 15

`define MRMAC__CTL_RX_MAX_PACKET_LEN_2    32'h000000df
`define MRMAC__CTL_RX_MAX_PACKET_LEN_2_SZ 15

`define MRMAC__CTL_RX_MAX_PACKET_LEN_3    32'h000000e0
`define MRMAC__CTL_RX_MAX_PACKET_LEN_3_SZ 15

`define MRMAC__CTL_RX_MIN_PACKET_LEN_0    32'h000000e1
`define MRMAC__CTL_RX_MIN_PACKET_LEN_0_SZ 8

`define MRMAC__CTL_RX_MIN_PACKET_LEN_1    32'h000000e2
`define MRMAC__CTL_RX_MIN_PACKET_LEN_1_SZ 8

`define MRMAC__CTL_RX_MIN_PACKET_LEN_2    32'h000000e3
`define MRMAC__CTL_RX_MIN_PACKET_LEN_2_SZ 8

`define MRMAC__CTL_RX_MIN_PACKET_LEN_3    32'h000000e4
`define MRMAC__CTL_RX_MIN_PACKET_LEN_3_SZ 8

`define MRMAC__CTL_RX_OPCODE_GPP_0    32'h000000e5
`define MRMAC__CTL_RX_OPCODE_GPP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_GPP_1    32'h000000e6
`define MRMAC__CTL_RX_OPCODE_GPP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_GPP_2    32'h000000e7
`define MRMAC__CTL_RX_OPCODE_GPP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_GPP_3    32'h000000e8
`define MRMAC__CTL_RX_OPCODE_GPP_3_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_GCP_0    32'h000000e9
`define MRMAC__CTL_RX_OPCODE_MAX_GCP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_GCP_1    32'h000000ea
`define MRMAC__CTL_RX_OPCODE_MAX_GCP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_GCP_2    32'h000000eb
`define MRMAC__CTL_RX_OPCODE_MAX_GCP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_GCP_3    32'h000000ec
`define MRMAC__CTL_RX_OPCODE_MAX_GCP_3_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_PCP_0    32'h000000ed
`define MRMAC__CTL_RX_OPCODE_MAX_PCP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_PCP_1    32'h000000ee
`define MRMAC__CTL_RX_OPCODE_MAX_PCP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_PCP_2    32'h000000ef
`define MRMAC__CTL_RX_OPCODE_MAX_PCP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_MAX_PCP_3    32'h000000f0
`define MRMAC__CTL_RX_OPCODE_MAX_PCP_3_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_GCP_0    32'h000000f1
`define MRMAC__CTL_RX_OPCODE_MIN_GCP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_GCP_1    32'h000000f2
`define MRMAC__CTL_RX_OPCODE_MIN_GCP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_GCP_2    32'h000000f3
`define MRMAC__CTL_RX_OPCODE_MIN_GCP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_GCP_3    32'h000000f4
`define MRMAC__CTL_RX_OPCODE_MIN_GCP_3_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_PCP_0    32'h000000f5
`define MRMAC__CTL_RX_OPCODE_MIN_PCP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_PCP_1    32'h000000f6
`define MRMAC__CTL_RX_OPCODE_MIN_PCP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_PCP_2    32'h000000f7
`define MRMAC__CTL_RX_OPCODE_MIN_PCP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_MIN_PCP_3    32'h000000f8
`define MRMAC__CTL_RX_OPCODE_MIN_PCP_3_SZ 16

`define MRMAC__CTL_RX_OPCODE_PPP_0    32'h000000f9
`define MRMAC__CTL_RX_OPCODE_PPP_0_SZ 16

`define MRMAC__CTL_RX_OPCODE_PPP_1    32'h000000fa
`define MRMAC__CTL_RX_OPCODE_PPP_1_SZ 16

`define MRMAC__CTL_RX_OPCODE_PPP_2    32'h000000fb
`define MRMAC__CTL_RX_OPCODE_PPP_2_SZ 16

`define MRMAC__CTL_RX_OPCODE_PPP_3    32'h000000fc
`define MRMAC__CTL_RX_OPCODE_PPP_3_SZ 16

`define MRMAC__CTL_RX_PAUSE_DA_MCAST_0    32'h000000fd
`define MRMAC__CTL_RX_PAUSE_DA_MCAST_0_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_MCAST_1    32'h000000fe
`define MRMAC__CTL_RX_PAUSE_DA_MCAST_1_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_MCAST_2    32'h000000ff
`define MRMAC__CTL_RX_PAUSE_DA_MCAST_2_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_MCAST_3    32'h00000100
`define MRMAC__CTL_RX_PAUSE_DA_MCAST_3_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_UCAST_0    32'h00000101
`define MRMAC__CTL_RX_PAUSE_DA_UCAST_0_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_UCAST_1    32'h00000102
`define MRMAC__CTL_RX_PAUSE_DA_UCAST_1_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_UCAST_2    32'h00000103
`define MRMAC__CTL_RX_PAUSE_DA_UCAST_2_SZ 48

`define MRMAC__CTL_RX_PAUSE_DA_UCAST_3    32'h00000104
`define MRMAC__CTL_RX_PAUSE_DA_UCAST_3_SZ 48

`define MRMAC__CTL_RX_PAUSE_SA_0    32'h00000105
`define MRMAC__CTL_RX_PAUSE_SA_0_SZ 48

`define MRMAC__CTL_RX_PAUSE_SA_1    32'h00000106
`define MRMAC__CTL_RX_PAUSE_SA_1_SZ 48

`define MRMAC__CTL_RX_PAUSE_SA_2    32'h00000107
`define MRMAC__CTL_RX_PAUSE_SA_2_SZ 48

`define MRMAC__CTL_RX_PAUSE_SA_3    32'h00000108
`define MRMAC__CTL_RX_PAUSE_SA_3_SZ 48

`define MRMAC__CTL_RX_PROCESS_LFI_0    32'h00000109
`define MRMAC__CTL_RX_PROCESS_LFI_0_SZ 40

`define MRMAC__CTL_RX_PROCESS_LFI_1    32'h0000010a
`define MRMAC__CTL_RX_PROCESS_LFI_1_SZ 40

`define MRMAC__CTL_RX_PROCESS_LFI_2    32'h0000010b
`define MRMAC__CTL_RX_PROCESS_LFI_2_SZ 40

`define MRMAC__CTL_RX_PROCESS_LFI_3    32'h0000010c
`define MRMAC__CTL_RX_PROCESS_LFI_3_SZ 40

`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_0    32'h0000010d
`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_0_SZ 20

`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_1    32'h0000010e
`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_1_SZ 20

`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_2    32'h0000010f
`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_2_SZ 20

`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_3    32'h00000110
`define MRMAC__CTL_RX_PTP_LATENCY_ADJUST_3_SZ 20

`define MRMAC__CTL_RX_PTP_ST_OFFSET_0    32'h00000111
`define MRMAC__CTL_RX_PTP_ST_OFFSET_0_SZ 16

`define MRMAC__CTL_RX_PTP_ST_OFFSET_1    32'h00000112
`define MRMAC__CTL_RX_PTP_ST_OFFSET_1_SZ 16

`define MRMAC__CTL_RX_PTP_ST_OFFSET_2    32'h00000113
`define MRMAC__CTL_RX_PTP_ST_OFFSET_2_SZ 16

`define MRMAC__CTL_RX_PTP_ST_OFFSET_3    32'h00000114
`define MRMAC__CTL_RX_PTP_ST_OFFSET_3_SZ 16

`define MRMAC__CTL_RX_TEST_PATTERN_0    32'h00000115
`define MRMAC__CTL_RX_TEST_PATTERN_0_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_1    32'h00000116
`define MRMAC__CTL_RX_TEST_PATTERN_1_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_2    32'h00000117
`define MRMAC__CTL_RX_TEST_PATTERN_2_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_3    32'h00000118
`define MRMAC__CTL_RX_TEST_PATTERN_3_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_0    32'h00000119
`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_0_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_1    32'h0000011a
`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_1_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_2    32'h0000011b
`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_2_SZ 40

`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_3    32'h0000011c
`define MRMAC__CTL_RX_TEST_PATTERN_ENABLE_3_SZ 40

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_100GE_0    32'h0000011d
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_100GE_0_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_0    32'h0000011e
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_0_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_1    32'h0000011f
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_1_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_2    32'h00000120
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_2_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_3    32'h00000121
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_25GE_3_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_40GE_0    32'h00000122
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_40GE_0_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_50GE_0    32'h00000123
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_50GE_0_SZ 16

`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_50GE_2    32'h00000124
`define MRMAC__CTL_RX_VL_LENGTH_MINUS1_50GE_2_SZ 16

`define MRMAC__CTL_SERDES_PASSTHRU_0    32'h00000125
`define MRMAC__CTL_SERDES_PASSTHRU_0_SZ 40

`define MRMAC__CTL_SERDES_PASSTHRU_1    32'h00000126
`define MRMAC__CTL_SERDES_PASSTHRU_1_SZ 40

`define MRMAC__CTL_SERDES_PASSTHRU_2    32'h00000127
`define MRMAC__CTL_SERDES_PASSTHRU_2_SZ 40

`define MRMAC__CTL_SERDES_PASSTHRU_3    32'h00000128
`define MRMAC__CTL_SERDES_PASSTHRU_3_SZ 40

`define MRMAC__CTL_SERDES_WIDTH_0    32'h00000129
`define MRMAC__CTL_SERDES_WIDTH_0_SZ 3

`define MRMAC__CTL_SERDES_WIDTH_1    32'h0000012a
`define MRMAC__CTL_SERDES_WIDTH_1_SZ 3

`define MRMAC__CTL_SERDES_WIDTH_2    32'h0000012b
`define MRMAC__CTL_SERDES_WIDTH_2_SZ 3

`define MRMAC__CTL_SERDES_WIDTH_3    32'h0000012c
`define MRMAC__CTL_SERDES_WIDTH_3_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_0    32'h0000012d
`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_0_SZ 4

`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_1    32'h0000012e
`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_1_SZ 4

`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_2    32'h0000012f
`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_2_SZ 4

`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_3    32'h00000130
`define MRMAC__CTL_TX_AXI_FIFO_HIGH_THRESHOLD_3_SZ 4

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_0    32'h00000131
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_0_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_1    32'h00000132
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_1_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_2    32'h00000133
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_2_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_3    32'h00000134
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_3_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_0    32'h00000135
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_0_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_1    32'h00000136
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_1_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_2    32'h00000137
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_2_SZ 3

`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_3    32'h00000138
`define MRMAC__CTL_TX_AXI_FIFO_LOW_THRESHOLD_ALT_3_SZ 3

`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_0    32'h00000139
`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_0_SZ 2

`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_1    32'h0000013a
`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_1_SZ 2

`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_2    32'h0000013b
`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_2_SZ 2

`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_3    32'h0000013c
`define MRMAC__CTL_TX_CORRUPT_FCS_ON_ERR_3_SZ 2

`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_0    32'h0000013d
`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_1    32'h0000013e
`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_2    32'h0000013f
`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_3    32'h00000140
`define MRMAC__CTL_TX_CUSTOM_PREAMBLE_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_0    32'h00000141
`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_0_SZ 40

`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_1    32'h00000142
`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_1_SZ 40

`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_2    32'h00000143
`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_2_SZ 40

`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_3    32'h00000144
`define MRMAC__CTL_TX_DATA_PATTERN_SELECT_3_SZ 40

`define MRMAC__CTL_TX_DA_GPP_0    32'h00000145
`define MRMAC__CTL_TX_DA_GPP_0_SZ 48

`define MRMAC__CTL_TX_DA_GPP_1    32'h00000146
`define MRMAC__CTL_TX_DA_GPP_1_SZ 48

`define MRMAC__CTL_TX_DA_GPP_2    32'h00000147
`define MRMAC__CTL_TX_DA_GPP_2_SZ 48

`define MRMAC__CTL_TX_DA_GPP_3    32'h00000148
`define MRMAC__CTL_TX_DA_GPP_3_SZ 48

`define MRMAC__CTL_TX_DA_PPP_0    32'h00000149
`define MRMAC__CTL_TX_DA_PPP_0_SZ 48

`define MRMAC__CTL_TX_DA_PPP_1    32'h0000014a
`define MRMAC__CTL_TX_DA_PPP_1_SZ 48

`define MRMAC__CTL_TX_DA_PPP_2    32'h0000014b
`define MRMAC__CTL_TX_DA_PPP_2_SZ 48

`define MRMAC__CTL_TX_DA_PPP_3    32'h0000014c
`define MRMAC__CTL_TX_DA_PPP_3_SZ 48

`define MRMAC__CTL_TX_ENABLE_0    32'h0000014d
`define MRMAC__CTL_TX_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_ENABLE_1    32'h0000014e
`define MRMAC__CTL_TX_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_ENABLE_2    32'h0000014f
`define MRMAC__CTL_TX_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_ENABLE_3    32'h00000150
`define MRMAC__CTL_TX_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_ETHERTYPE_GPP_0    32'h00000151
`define MRMAC__CTL_TX_ETHERTYPE_GPP_0_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_GPP_1    32'h00000152
`define MRMAC__CTL_TX_ETHERTYPE_GPP_1_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_GPP_2    32'h00000153
`define MRMAC__CTL_TX_ETHERTYPE_GPP_2_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_GPP_3    32'h00000154
`define MRMAC__CTL_TX_ETHERTYPE_GPP_3_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_PPP_0    32'h00000155
`define MRMAC__CTL_TX_ETHERTYPE_PPP_0_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_PPP_1    32'h00000156
`define MRMAC__CTL_TX_ETHERTYPE_PPP_1_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_PPP_2    32'h00000157
`define MRMAC__CTL_TX_ETHERTYPE_PPP_2_SZ 16

`define MRMAC__CTL_TX_ETHERTYPE_PPP_3    32'h00000158
`define MRMAC__CTL_TX_ETHERTYPE_PPP_3_SZ 16

`define MRMAC__CTL_TX_FCS_INS_ENABLE_0    32'h00000159
`define MRMAC__CTL_TX_FCS_INS_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_FCS_INS_ENABLE_1    32'h0000015a
`define MRMAC__CTL_TX_FCS_INS_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_FCS_INS_ENABLE_2    32'h0000015b
`define MRMAC__CTL_TX_FCS_INS_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_FCS_INS_ENABLE_3    32'h0000015c
`define MRMAC__CTL_TX_FCS_INS_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_FEC_FOUR_LANE_PMD    32'h0000015d
`define MRMAC__CTL_TX_FEC_FOUR_LANE_PMD_SZ 40

`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_0    32'h0000015e
`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_0_SZ 40

`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_1    32'h0000015f
`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_1_SZ 40

`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_2    32'h00000160
`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_2_SZ 40

`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_3    32'h00000161
`define MRMAC__CTL_TX_FEC_TRANSCODE_BYPASS_3_SZ 40

`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_0    32'h00000162
`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_1    32'h00000163
`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_2    32'h00000164
`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_3    32'h00000165
`define MRMAC__CTL_TX_FLEXIF_INPUT_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_FLEXIF_SELECT_0    32'h00000166
`define MRMAC__CTL_TX_FLEXIF_SELECT_0_SZ 3

`define MRMAC__CTL_TX_FLEXIF_SELECT_1    32'h00000167
`define MRMAC__CTL_TX_FLEXIF_SELECT_1_SZ 3

`define MRMAC__CTL_TX_FLEXIF_SELECT_2    32'h00000168
`define MRMAC__CTL_TX_FLEXIF_SELECT_2_SZ 3

`define MRMAC__CTL_TX_FLEXIF_SELECT_3    32'h00000169
`define MRMAC__CTL_TX_FLEXIF_SELECT_3_SZ 3

`define MRMAC__CTL_TX_IGNORE_FCS_0    32'h0000016a
`define MRMAC__CTL_TX_IGNORE_FCS_0_SZ 40

`define MRMAC__CTL_TX_IGNORE_FCS_1    32'h0000016b
`define MRMAC__CTL_TX_IGNORE_FCS_1_SZ 40

`define MRMAC__CTL_TX_IGNORE_FCS_2    32'h0000016c
`define MRMAC__CTL_TX_IGNORE_FCS_2_SZ 40

`define MRMAC__CTL_TX_IGNORE_FCS_3    32'h0000016d
`define MRMAC__CTL_TX_IGNORE_FCS_3_SZ 40

`define MRMAC__CTL_TX_IPG_VALUE_0    32'h0000016e
`define MRMAC__CTL_TX_IPG_VALUE_0_SZ 4

`define MRMAC__CTL_TX_IPG_VALUE_1    32'h0000016f
`define MRMAC__CTL_TX_IPG_VALUE_1_SZ 4

`define MRMAC__CTL_TX_IPG_VALUE_2    32'h00000170
`define MRMAC__CTL_TX_IPG_VALUE_2_SZ 4

`define MRMAC__CTL_TX_IPG_VALUE_3    32'h00000171
`define MRMAC__CTL_TX_IPG_VALUE_3_SZ 4

`define MRMAC__CTL_TX_OPCODE_GPP_0    32'h00000172
`define MRMAC__CTL_TX_OPCODE_GPP_0_SZ 16

`define MRMAC__CTL_TX_OPCODE_GPP_1    32'h00000173
`define MRMAC__CTL_TX_OPCODE_GPP_1_SZ 16

`define MRMAC__CTL_TX_OPCODE_GPP_2    32'h00000174
`define MRMAC__CTL_TX_OPCODE_GPP_2_SZ 16

`define MRMAC__CTL_TX_OPCODE_GPP_3    32'h00000175
`define MRMAC__CTL_TX_OPCODE_GPP_3_SZ 16

`define MRMAC__CTL_TX_OPCODE_PPP_0    32'h00000176
`define MRMAC__CTL_TX_OPCODE_PPP_0_SZ 16

`define MRMAC__CTL_TX_OPCODE_PPP_1    32'h00000177
`define MRMAC__CTL_TX_OPCODE_PPP_1_SZ 16

`define MRMAC__CTL_TX_OPCODE_PPP_2    32'h00000178
`define MRMAC__CTL_TX_OPCODE_PPP_2_SZ 16

`define MRMAC__CTL_TX_OPCODE_PPP_3    32'h00000179
`define MRMAC__CTL_TX_OPCODE_PPP_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA0_0    32'h0000017a
`define MRMAC__CTL_TX_PAUSE_QUANTA0_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA0_1    32'h0000017b
`define MRMAC__CTL_TX_PAUSE_QUANTA0_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA0_2    32'h0000017c
`define MRMAC__CTL_TX_PAUSE_QUANTA0_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA0_3    32'h0000017d
`define MRMAC__CTL_TX_PAUSE_QUANTA0_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA1_0    32'h0000017e
`define MRMAC__CTL_TX_PAUSE_QUANTA1_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA1_1    32'h0000017f
`define MRMAC__CTL_TX_PAUSE_QUANTA1_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA1_2    32'h00000180
`define MRMAC__CTL_TX_PAUSE_QUANTA1_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA1_3    32'h00000181
`define MRMAC__CTL_TX_PAUSE_QUANTA1_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA2_0    32'h00000182
`define MRMAC__CTL_TX_PAUSE_QUANTA2_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA2_1    32'h00000183
`define MRMAC__CTL_TX_PAUSE_QUANTA2_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA2_2    32'h00000184
`define MRMAC__CTL_TX_PAUSE_QUANTA2_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA2_3    32'h00000185
`define MRMAC__CTL_TX_PAUSE_QUANTA2_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA3_0    32'h00000186
`define MRMAC__CTL_TX_PAUSE_QUANTA3_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA3_1    32'h00000187
`define MRMAC__CTL_TX_PAUSE_QUANTA3_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA3_2    32'h00000188
`define MRMAC__CTL_TX_PAUSE_QUANTA3_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA3_3    32'h00000189
`define MRMAC__CTL_TX_PAUSE_QUANTA3_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA4_0    32'h0000018a
`define MRMAC__CTL_TX_PAUSE_QUANTA4_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA4_1    32'h0000018b
`define MRMAC__CTL_TX_PAUSE_QUANTA4_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA4_2    32'h0000018c
`define MRMAC__CTL_TX_PAUSE_QUANTA4_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA4_3    32'h0000018d
`define MRMAC__CTL_TX_PAUSE_QUANTA4_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA5_0    32'h0000018e
`define MRMAC__CTL_TX_PAUSE_QUANTA5_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA5_1    32'h0000018f
`define MRMAC__CTL_TX_PAUSE_QUANTA5_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA5_2    32'h00000190
`define MRMAC__CTL_TX_PAUSE_QUANTA5_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA5_3    32'h00000191
`define MRMAC__CTL_TX_PAUSE_QUANTA5_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA6_0    32'h00000192
`define MRMAC__CTL_TX_PAUSE_QUANTA6_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA6_1    32'h00000193
`define MRMAC__CTL_TX_PAUSE_QUANTA6_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA6_2    32'h00000194
`define MRMAC__CTL_TX_PAUSE_QUANTA6_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA6_3    32'h00000195
`define MRMAC__CTL_TX_PAUSE_QUANTA6_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA7_0    32'h00000196
`define MRMAC__CTL_TX_PAUSE_QUANTA7_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA7_1    32'h00000197
`define MRMAC__CTL_TX_PAUSE_QUANTA7_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA7_2    32'h00000198
`define MRMAC__CTL_TX_PAUSE_QUANTA7_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA7_3    32'h00000199
`define MRMAC__CTL_TX_PAUSE_QUANTA7_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA8_0    32'h0000019a
`define MRMAC__CTL_TX_PAUSE_QUANTA8_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA8_1    32'h0000019b
`define MRMAC__CTL_TX_PAUSE_QUANTA8_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA8_2    32'h0000019c
`define MRMAC__CTL_TX_PAUSE_QUANTA8_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_QUANTA8_3    32'h0000019d
`define MRMAC__CTL_TX_PAUSE_QUANTA8_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_0    32'h0000019e
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_1    32'h0000019f
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_2    32'h000001a0
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_3    32'h000001a1
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER0_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_0    32'h000001a2
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_1    32'h000001a3
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_2    32'h000001a4
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_3    32'h000001a5
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER1_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_0    32'h000001a6
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_1    32'h000001a7
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_2    32'h000001a8
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_3    32'h000001a9
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER2_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_0    32'h000001aa
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_1    32'h000001ab
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_2    32'h000001ac
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_3    32'h000001ad
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER3_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_0    32'h000001ae
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_1    32'h000001af
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_2    32'h000001b0
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_3    32'h000001b1
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER4_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_0    32'h000001b2
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_1    32'h000001b3
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_2    32'h000001b4
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_3    32'h000001b5
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER5_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_0    32'h000001b6
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_1    32'h000001b7
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_2    32'h000001b8
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_3    32'h000001b9
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER6_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_0    32'h000001ba
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_1    32'h000001bb
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_2    32'h000001bc
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_3    32'h000001bd
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER7_3_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_0    32'h000001be
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_0_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_1    32'h000001bf
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_1_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_2    32'h000001c0
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_2_SZ 16

`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_3    32'h000001c1
`define MRMAC__CTL_TX_PAUSE_REFRESH_TIMER8_3_SZ 16

`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_0    32'h000001c2
`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_1    32'h000001c3
`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_2    32'h000001c4
`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_3    32'h000001c5
`define MRMAC__CTL_TX_PTP_1STEP_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_0    32'h000001c6
`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_0_SZ 20

`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_1    32'h000001c7
`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_1_SZ 20

`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_2    32'h000001c8
`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_2_SZ 20

`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_3    32'h000001c9
`define MRMAC__CTL_TX_PTP_LATENCY_ADJUST_3_SZ 20

`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_0    32'h000001ca
`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_0_SZ 40

`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_1    32'h000001cb
`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_1_SZ 40

`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_2    32'h000001cc
`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_2_SZ 40

`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_3    32'h000001cd
`define MRMAC__CTL_TX_PTP_RSFEC_COMP_EN_3_SZ 40

`define MRMAC__CTL_TX_PTP_SAT_ENABLE_0    32'h000001ce
`define MRMAC__CTL_TX_PTP_SAT_ENABLE_0_SZ 2

`define MRMAC__CTL_TX_PTP_SAT_ENABLE_1    32'h000001cf
`define MRMAC__CTL_TX_PTP_SAT_ENABLE_1_SZ 2

`define MRMAC__CTL_TX_PTP_SAT_ENABLE_2    32'h000001d0
`define MRMAC__CTL_TX_PTP_SAT_ENABLE_2_SZ 2

`define MRMAC__CTL_TX_PTP_SAT_ENABLE_3    32'h000001d1
`define MRMAC__CTL_TX_PTP_SAT_ENABLE_3_SZ 2

`define MRMAC__CTL_TX_PTP_ST_OFFSET_0    32'h000001d2
`define MRMAC__CTL_TX_PTP_ST_OFFSET_0_SZ 16

`define MRMAC__CTL_TX_PTP_ST_OFFSET_1    32'h000001d3
`define MRMAC__CTL_TX_PTP_ST_OFFSET_1_SZ 16

`define MRMAC__CTL_TX_PTP_ST_OFFSET_2    32'h000001d4
`define MRMAC__CTL_TX_PTP_ST_OFFSET_2_SZ 16

`define MRMAC__CTL_TX_PTP_ST_OFFSET_3    32'h000001d5
`define MRMAC__CTL_TX_PTP_ST_OFFSET_3_SZ 16

`define MRMAC__CTL_TX_SA_GPP_0    32'h000001d6
`define MRMAC__CTL_TX_SA_GPP_0_SZ 48

`define MRMAC__CTL_TX_SA_GPP_1    32'h000001d7
`define MRMAC__CTL_TX_SA_GPP_1_SZ 48

`define MRMAC__CTL_TX_SA_GPP_2    32'h000001d8
`define MRMAC__CTL_TX_SA_GPP_2_SZ 48

`define MRMAC__CTL_TX_SA_GPP_3    32'h000001d9
`define MRMAC__CTL_TX_SA_GPP_3_SZ 48

`define MRMAC__CTL_TX_SA_PPP_0    32'h000001da
`define MRMAC__CTL_TX_SA_PPP_0_SZ 48

`define MRMAC__CTL_TX_SA_PPP_1    32'h000001db
`define MRMAC__CTL_TX_SA_PPP_1_SZ 48

`define MRMAC__CTL_TX_SA_PPP_2    32'h000001dc
`define MRMAC__CTL_TX_SA_PPP_2_SZ 48

`define MRMAC__CTL_TX_SA_PPP_3    32'h000001dd
`define MRMAC__CTL_TX_SA_PPP_3_SZ 48

`define MRMAC__CTL_TX_SEND_IDLE_0    32'h000001de
`define MRMAC__CTL_TX_SEND_IDLE_0_SZ 40

`define MRMAC__CTL_TX_SEND_IDLE_1    32'h000001df
`define MRMAC__CTL_TX_SEND_IDLE_1_SZ 40

`define MRMAC__CTL_TX_SEND_IDLE_2    32'h000001e0
`define MRMAC__CTL_TX_SEND_IDLE_2_SZ 40

`define MRMAC__CTL_TX_SEND_IDLE_3    32'h000001e1
`define MRMAC__CTL_TX_SEND_IDLE_3_SZ 40

`define MRMAC__CTL_TX_SEND_LFI_0    32'h000001e2
`define MRMAC__CTL_TX_SEND_LFI_0_SZ 40

`define MRMAC__CTL_TX_SEND_LFI_1    32'h000001e3
`define MRMAC__CTL_TX_SEND_LFI_1_SZ 40

`define MRMAC__CTL_TX_SEND_LFI_2    32'h000001e4
`define MRMAC__CTL_TX_SEND_LFI_2_SZ 40

`define MRMAC__CTL_TX_SEND_LFI_3    32'h000001e5
`define MRMAC__CTL_TX_SEND_LFI_3_SZ 40

`define MRMAC__CTL_TX_SEND_RFI_0    32'h000001e6
`define MRMAC__CTL_TX_SEND_RFI_0_SZ 40

`define MRMAC__CTL_TX_SEND_RFI_1    32'h000001e7
`define MRMAC__CTL_TX_SEND_RFI_1_SZ 40

`define MRMAC__CTL_TX_SEND_RFI_2    32'h000001e8
`define MRMAC__CTL_TX_SEND_RFI_2_SZ 40

`define MRMAC__CTL_TX_SEND_RFI_3    32'h000001e9
`define MRMAC__CTL_TX_SEND_RFI_3_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_0    32'h000001ea
`define MRMAC__CTL_TX_TEST_PATTERN_0_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_1    32'h000001eb
`define MRMAC__CTL_TX_TEST_PATTERN_1_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_2    32'h000001ec
`define MRMAC__CTL_TX_TEST_PATTERN_2_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_3    32'h000001ed
`define MRMAC__CTL_TX_TEST_PATTERN_3_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_0    32'h000001ee
`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_0_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_1    32'h000001ef
`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_1_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_2    32'h000001f0
`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_2_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_3    32'h000001f1
`define MRMAC__CTL_TX_TEST_PATTERN_ENABLE_3_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_0    32'h000001f2
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_0_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_1    32'h000001f3
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_1_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_2    32'h000001f4
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_2_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_3    32'h000001f5
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_A_3_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_0    32'h000001f6
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_0_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_1    32'h000001f7
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_1_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_2    32'h000001f8
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_2_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_3    32'h000001f9
`define MRMAC__CTL_TX_TEST_PATTERN_SEED_B_3_SZ 58

`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_0    32'h000001fa
`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_0_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_1    32'h000001fb
`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_1_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_2    32'h000001fc
`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_2_SZ 40

`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_3    32'h000001fd
`define MRMAC__CTL_TX_TEST_PATTERN_SELECT_3_SZ 40

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_100GE_0    32'h000001fe
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_100GE_0_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_0    32'h000001ff
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_0_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_1    32'h00000200
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_1_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_2    32'h00000201
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_2_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_3    32'h00000202
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_25GE_3_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_40GE_0    32'h00000203
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_40GE_0_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_50GE_0    32'h00000204
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_50GE_0_SZ 16

`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_50GE_2    32'h00000205
`define MRMAC__CTL_TX_VL_LENGTH_MINUS1_50GE_2_SZ 16

`define MRMAC__CTL_VL_MARKER_ID0    32'h00000206
`define MRMAC__CTL_VL_MARKER_ID0_SZ 64

`define MRMAC__CTL_VL_MARKER_ID1    32'h00000207
`define MRMAC__CTL_VL_MARKER_ID1_SZ 64

`define MRMAC__CTL_VL_MARKER_ID10    32'h00000208
`define MRMAC__CTL_VL_MARKER_ID10_SZ 64

`define MRMAC__CTL_VL_MARKER_ID11    32'h00000209
`define MRMAC__CTL_VL_MARKER_ID11_SZ 64

`define MRMAC__CTL_VL_MARKER_ID12    32'h0000020a
`define MRMAC__CTL_VL_MARKER_ID12_SZ 64

`define MRMAC__CTL_VL_MARKER_ID13    32'h0000020b
`define MRMAC__CTL_VL_MARKER_ID13_SZ 64

`define MRMAC__CTL_VL_MARKER_ID14    32'h0000020c
`define MRMAC__CTL_VL_MARKER_ID14_SZ 64

`define MRMAC__CTL_VL_MARKER_ID15    32'h0000020d
`define MRMAC__CTL_VL_MARKER_ID15_SZ 64

`define MRMAC__CTL_VL_MARKER_ID16    32'h0000020e
`define MRMAC__CTL_VL_MARKER_ID16_SZ 64

`define MRMAC__CTL_VL_MARKER_ID17    32'h0000020f
`define MRMAC__CTL_VL_MARKER_ID17_SZ 64

`define MRMAC__CTL_VL_MARKER_ID18    32'h00000210
`define MRMAC__CTL_VL_MARKER_ID18_SZ 64

`define MRMAC__CTL_VL_MARKER_ID19    32'h00000211
`define MRMAC__CTL_VL_MARKER_ID19_SZ 64

`define MRMAC__CTL_VL_MARKER_ID2    32'h00000212
`define MRMAC__CTL_VL_MARKER_ID2_SZ 64

`define MRMAC__CTL_VL_MARKER_ID3    32'h00000213
`define MRMAC__CTL_VL_MARKER_ID3_SZ 64

`define MRMAC__CTL_VL_MARKER_ID4    32'h00000214
`define MRMAC__CTL_VL_MARKER_ID4_SZ 64

`define MRMAC__CTL_VL_MARKER_ID5    32'h00000215
`define MRMAC__CTL_VL_MARKER_ID5_SZ 64

`define MRMAC__CTL_VL_MARKER_ID6    32'h00000216
`define MRMAC__CTL_VL_MARKER_ID6_SZ 64

`define MRMAC__CTL_VL_MARKER_ID7    32'h00000217
`define MRMAC__CTL_VL_MARKER_ID7_SZ 64

`define MRMAC__CTL_VL_MARKER_ID8    32'h00000218
`define MRMAC__CTL_VL_MARKER_ID8_SZ 64

`define MRMAC__CTL_VL_MARKER_ID9    32'h00000219
`define MRMAC__CTL_VL_MARKER_ID9_SZ 64

`define MRMAC__LANE_CONNECTIVITY    32'h0000021a
`define MRMAC__LANE_CONNECTIVITY_SZ 32

`define MRMAC__MEM_CTRL    32'h0000021b
`define MRMAC__MEM_CTRL_SZ 8

`define MRMAC__NUM_100G_FEC_ONLY_PORTS    32'h0000021c
`define MRMAC__NUM_100G_FEC_ONLY_PORTS_SZ 1

`define MRMAC__NUM_100G_MAC_PCS_NOFEC_PORTS    32'h0000021d
`define MRMAC__NUM_100G_MAC_PCS_NOFEC_PORTS_SZ 1

`define MRMAC__NUM_100G_MAC_PCS_WITH_FEC_PORTS    32'h0000021e
`define MRMAC__NUM_100G_MAC_PCS_WITH_FEC_PORTS_SZ 1

`define MRMAC__NUM_10G_MAC_PCS_NOFEC_PORTS    32'h0000021f
`define MRMAC__NUM_10G_MAC_PCS_NOFEC_PORTS_SZ 3

`define MRMAC__NUM_10G_MAC_PCS_WITH_FEC_PORTS    32'h00000220
`define MRMAC__NUM_10G_MAC_PCS_WITH_FEC_PORTS_SZ 3

`define MRMAC__NUM_25G_FEC_ONLY_PORTS    32'h00000221
`define MRMAC__NUM_25G_FEC_ONLY_PORTS_SZ 3

`define MRMAC__NUM_25G_MAC_PCS_NOFEC_PORTS    32'h00000222
`define MRMAC__NUM_25G_MAC_PCS_NOFEC_PORTS_SZ 3

`define MRMAC__NUM_25G_MAC_PCS_WITH_FEC_PORTS    32'h00000223
`define MRMAC__NUM_25G_MAC_PCS_WITH_FEC_PORTS_SZ 3

`define MRMAC__NUM_40G_MAC_PCS_NOFEC_PORTS    32'h00000224
`define MRMAC__NUM_40G_MAC_PCS_NOFEC_PORTS_SZ 1

`define MRMAC__NUM_40G_MAC_PCS_WITH_FEC_PORTS    32'h00000225
`define MRMAC__NUM_40G_MAC_PCS_WITH_FEC_PORTS_SZ 1

`define MRMAC__NUM_50G_FEC_ONLY_PORTS    32'h00000226
`define MRMAC__NUM_50G_FEC_ONLY_PORTS_SZ 2

`define MRMAC__NUM_50G_MAC_PCS_NOFEC_PORTS    32'h00000227
`define MRMAC__NUM_50G_MAC_PCS_NOFEC_PORTS_SZ 2

`define MRMAC__NUM_50G_MAC_PCS_WITH_FEC_PORTS    32'h00000228
`define MRMAC__NUM_50G_MAC_PCS_WITH_FEC_PORTS_SZ 2

`define MRMAC__RSVD0    32'h00000229
`define MRMAC__RSVD0_SZ 32

`define MRMAC__RSVD1    32'h0000022a
`define MRMAC__RSVD1_SZ 32

`define MRMAC__RSVD2    32'h0000022b
`define MRMAC__RSVD2_SZ 32

`define MRMAC__RSVD3    32'h0000022c
`define MRMAC__RSVD3_SZ 32

`define MRMAC__RSVD4    32'h0000022d
`define MRMAC__RSVD4_SZ 32

`define MRMAC__RSVD5    32'h0000022e
`define MRMAC__RSVD5_SZ 32

`define MRMAC__RSVD6    32'h0000022f
`define MRMAC__RSVD6_SZ 32

`define MRMAC__RSVD7    32'h00000230
`define MRMAC__RSVD7_SZ 32

`define MRMAC__RSVD8    32'h00000231
`define MRMAC__RSVD8_SZ 32

`define MRMAC__RSVD9    32'h00000232
`define MRMAC__RSVD9_SZ 32

`define MRMAC__SIM_DEVICE    32'h00000233
`define MRMAC__SIM_DEVICE_SZ 144

`define MRMAC__TICK_REG_MODE_SEL_0    32'h00000234
`define MRMAC__TICK_REG_MODE_SEL_0_SZ 40

`define MRMAC__TICK_REG_MODE_SEL_1    32'h00000235
`define MRMAC__TICK_REG_MODE_SEL_1_SZ 40

`define MRMAC__TICK_REG_MODE_SEL_2    32'h00000236
`define MRMAC__TICK_REG_MODE_SEL_2_SZ 40

`define MRMAC__TICK_REG_MODE_SEL_3    32'h00000237
`define MRMAC__TICK_REG_MODE_SEL_3_SZ 40

`endif  // B_MRMAC_DEFINES_VH