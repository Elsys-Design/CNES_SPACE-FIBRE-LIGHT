----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/03/2024
--
-- Description : This module compute the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

entity data_seq_compute is
port (
	RST_N                 : in  std_logic;                                    --! global reset
	CLK                   : in  std_logic;                                    --! Clock generated by GTY IP
	-- Lane Interface
	LANE_ACTIVE_PPL       : in  std_logic;                                    --! Lane Active flag for the DATA Link Layer
	-- DENC interface
	NEW_WORD_DENC         : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
	DATA_DENC             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
	VALID_K_CHARAC_DENC   : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
	TYPE_FRAME_DENC       : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
	END_FRAME_DENC        : in  std_logic;
	-- DENC interface
	NEW_WORD_DSCOM        : out  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
	DATA_DSCOM            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
	VALID_K_CHARAC_DSCOM  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
	TYPE_FRAME_DSCOM      : out  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
	END_FRAME_DSCOM       : out  std_logic;
	-- MIB interface
	SEQ_NUM_DSCOM         : out std_logic_vector(7 downto 0)
  );
end data_seq_compute;

architecture rtl of data_seq_compute is
---------------------------------------------------------
-----                  Declaration signals          -----
---------------------------------------------------------

signal trans_seq_cnt    : unsigned(6 downto 0);   --! Data parallel from Lane Layer
signal trans_pol_flg    : std_logic;               --! Data parallel from Lane Layer
begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_seq_num_comp
-- Description: Comute the SEQ_NUM for each frame
---------------------------------------------------------
p_seq_num_comp: process(CLK, RST_N)
begin
	if RST_N = '0' then
	  trans_seq_cnt        <= (others => '0'); -- Reset seq_num_cnt	on link reset
		trans_pol_flg        <= '0';
		NEW_WORD_DSCOM       <= '0';
		VALID_K_CHARAC_DSCOM <= (others => '0');
		TYPE_FRAME_DSCOM     <= (others => '0');
		END_FRAME_DSCOM      <= '0';
		DATA_DSCOM           <= (others => '0');
		SEQ_NUM_DSCOM        <= (others => '0');
	elsif rising_edge(CLK) and LANE_ACTIVE_PPL= '1' then
		NEW_WORD_DSCOM       <= NEW_WORD_DENC;
		VALID_K_CHARAC_DSCOM <= VALID_K_CHARAC_DENC;
		TYPE_FRAME_DSCOM     <= TYPE_FRAME_DENC;
		END_FRAME_DSCOM      <= END_FRAME_DENC;
		if END_FRAME_DENC = '1' then -- control word or EDF or EBF
			if TYPE_FRAME_DENC = C_DATA_FRM then
				DATA_DSCOM      <= C_RESERVED_SYMB & C_RESERVED_SYMB & trans_pol_flg & std_logic_vector(trans_seq_cnt+1) & DATA_DENC(7 downto 0);
				SEQ_NUM_DSCOM   <= trans_pol_flg & std_logic_vector(trans_seq_cnt+1);
				trans_seq_cnt   <= trans_seq_cnt +1;
			elsif TYPE_FRAME_DENC = C_BC_FRM or TYPE_FRAME_DENC = C_FCT_FRM then
				DATA_DSCOM      <= C_RESERVED_SYMB & trans_pol_flg & std_logic_vector(trans_seq_cnt+1) & DATA_DENC(15 downto 0);
				SEQ_NUM_DSCOM   <= trans_pol_flg & std_logic_vector(trans_seq_cnt+1);
				trans_seq_cnt   <= trans_seq_cnt +1;
			else
				DATA_DSCOM      <= C_RESERVED_SYMB & trans_pol_flg & std_logic_vector(trans_seq_cnt) & DATA_DENC(15 downto 0);
				SEQ_NUM_DSCOM   <= trans_pol_flg & std_logic_vector(trans_seq_cnt);
			end if;
		elsif DATA_DENC(7 downto 0) = C_K28_7_SYMB and VALID_K_CHARAC_DENC(0)= '1' then -- SIF or SDF or SBF
			DATA_DSCOM      <= C_RESERVED_SYMB & trans_pol_flg & std_logic_vector(trans_seq_cnt) & DATA_DENC(15 downto 0);
			SEQ_NUM_DSCOM   <= trans_pol_flg & std_logic_vector(trans_seq_cnt);
		else
      DATA_DSCOM      <= DATA_DENC;
		end if;
	end if;
end process p_seq_num_comp;

end architecture rtl;