`include "B_HBM_SNGLBLI_INTF_APB_defines.vh"

reg [`HBM_SNGLBLI_INTF_APB_DATA_SZ-1:0] ATTR [0:`HBM_SNGLBLI_INTF_APB_ADDR_N-1];
reg [`HBM_SNGLBLI_INTF_APB__CLK_SEL_SZ:1] CLK_SEL_REG = CLK_SEL;
reg IS_PCLK_INVERTED_REG = IS_PCLK_INVERTED;
reg IS_PRESET_N_INVERTED_REG = IS_PRESET_N_INVERTED;
reg [`HBM_SNGLBLI_INTF_APB__MC_ENABLE_SZ:1] MC_ENABLE_REG = MC_ENABLE;
reg [`HBM_SNGLBLI_INTF_APB__PHY_ENABLE_SZ:1] PHY_ENABLE_REG = PHY_ENABLE;
reg [`HBM_SNGLBLI_INTF_APB__PHY_PCLK_INVERT_SZ:1] PHY_PCLK_INVERT_REG = PHY_PCLK_INVERT;
reg [`HBM_SNGLBLI_INTF_APB__SWITCH_ENABLE_SZ:1] SWITCH_ENABLE_REG = SWITCH_ENABLE;

initial begin
  ATTR[`HBM_SNGLBLI_INTF_APB__CLK_SEL] = CLK_SEL;
  ATTR[`HBM_SNGLBLI_INTF_APB__IS_PCLK_INVERTED] = IS_PCLK_INVERTED;
  ATTR[`HBM_SNGLBLI_INTF_APB__IS_PRESET_N_INVERTED] = IS_PRESET_N_INVERTED;
  ATTR[`HBM_SNGLBLI_INTF_APB__MC_ENABLE] = MC_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_APB__PHY_ENABLE] = PHY_ENABLE;
  ATTR[`HBM_SNGLBLI_INTF_APB__PHY_PCLK_INVERT] = PHY_PCLK_INVERT;
  ATTR[`HBM_SNGLBLI_INTF_APB__SWITCH_ENABLE] = SWITCH_ENABLE;
end

always @(trig_attr) begin
  CLK_SEL_REG = ATTR[`HBM_SNGLBLI_INTF_APB__CLK_SEL];
  IS_PCLK_INVERTED_REG = ATTR[`HBM_SNGLBLI_INTF_APB__IS_PCLK_INVERTED];
  IS_PRESET_N_INVERTED_REG = ATTR[`HBM_SNGLBLI_INTF_APB__IS_PRESET_N_INVERTED];
  MC_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_APB__MC_ENABLE];
  PHY_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_APB__PHY_ENABLE];
  PHY_PCLK_INVERT_REG = ATTR[`HBM_SNGLBLI_INTF_APB__PHY_PCLK_INVERT];
  SWITCH_ENABLE_REG = ATTR[`HBM_SNGLBLI_INTF_APB__SWITCH_ENABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`HBM_SNGLBLI_INTF_APB_ADDR_SZ-1:0] addr;
  input  [`HBM_SNGLBLI_INTF_APB_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`HBM_SNGLBLI_INTF_APB_DATA_SZ-1:0] read_attr;
  input  [`HBM_SNGLBLI_INTF_APB_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
