`include "B_ODELAYE2_defines.vh"

reg [`ODELAYE2_DATA_SZ-1:0] ATTR [0:`ODELAYE2_ADDR_N-1];
reg [`ODELAYE2__CINVCTRL_SEL_SZ:1] CINVCTRL_SEL_REG = CINVCTRL_SEL;
reg [`ODELAYE2__DELAY_SRC_SZ:1] DELAY_SRC_REG = DELAY_SRC;
reg [`ODELAYE2__HIGH_PERFORMANCE_MODE_SZ:1] HIGH_PERFORMANCE_MODE_REG = HIGH_PERFORMANCE_MODE;
reg IS_C_INVERTED_REG = IS_C_INVERTED;
reg IS_ODATAIN_INVERTED_REG = IS_ODATAIN_INVERTED;
reg [`ODELAYE2__ODELAY_TYPE_SZ:1] ODELAY_TYPE_REG = ODELAY_TYPE;
reg [`ODELAYE2__ODELAY_VALUE_SZ-1:0] ODELAY_VALUE_REG = ODELAY_VALUE;
reg [`ODELAYE2__PIPE_SEL_SZ:1] PIPE_SEL_REG = PIPE_SEL;
real REFCLK_FREQUENCY_REG = REFCLK_FREQUENCY;
reg [`ODELAYE2__SIGNAL_PATTERN_SZ:1] SIGNAL_PATTERN_REG = SIGNAL_PATTERN;
reg [`ODELAYE2__SIM_DELAY_D_SZ-1:0] SIM_DELAY_D_REG = SIM_DELAY_D;

initial begin
  ATTR[`ODELAYE2__CINVCTRL_SEL] = CINVCTRL_SEL;
  ATTR[`ODELAYE2__DELAY_SRC] = DELAY_SRC;
  ATTR[`ODELAYE2__HIGH_PERFORMANCE_MODE] = HIGH_PERFORMANCE_MODE;
  ATTR[`ODELAYE2__IS_C_INVERTED] = IS_C_INVERTED;
  ATTR[`ODELAYE2__IS_ODATAIN_INVERTED] = IS_ODATAIN_INVERTED;
  ATTR[`ODELAYE2__ODELAY_TYPE] = ODELAY_TYPE;
  ATTR[`ODELAYE2__ODELAY_VALUE] = ODELAY_VALUE;
  ATTR[`ODELAYE2__PIPE_SEL] = PIPE_SEL;
  ATTR[`ODELAYE2__REFCLK_FREQUENCY] = $realtobits(REFCLK_FREQUENCY);
  ATTR[`ODELAYE2__SIGNAL_PATTERN] = SIGNAL_PATTERN;
  ATTR[`ODELAYE2__SIM_DELAY_D] = SIM_DELAY_D;
end

always @(trig_attr) begin
  CINVCTRL_SEL_REG = ATTR[`ODELAYE2__CINVCTRL_SEL];
  DELAY_SRC_REG = ATTR[`ODELAYE2__DELAY_SRC];
  HIGH_PERFORMANCE_MODE_REG = ATTR[`ODELAYE2__HIGH_PERFORMANCE_MODE];
  IS_C_INVERTED_REG = ATTR[`ODELAYE2__IS_C_INVERTED];
  IS_ODATAIN_INVERTED_REG = ATTR[`ODELAYE2__IS_ODATAIN_INVERTED];
  ODELAY_TYPE_REG = ATTR[`ODELAYE2__ODELAY_TYPE];
  ODELAY_VALUE_REG = ATTR[`ODELAYE2__ODELAY_VALUE];
  PIPE_SEL_REG = ATTR[`ODELAYE2__PIPE_SEL];
  REFCLK_FREQUENCY_REG = $bitstoreal(ATTR[`ODELAYE2__REFCLK_FREQUENCY]);
  SIGNAL_PATTERN_REG = ATTR[`ODELAYE2__SIGNAL_PATTERN];
  SIM_DELAY_D_REG = ATTR[`ODELAYE2__SIM_DELAY_D];
end

// procedures to override, read attribute values

task write_attr;
  input  [`ODELAYE2_ADDR_SZ-1:0] addr;
  input  [`ODELAYE2_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`ODELAYE2_DATA_SZ-1:0] read_attr;
  input  [`ODELAYE2_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
