// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP58_DEFINES_VH
`else
`define B_DSP58_DEFINES_VH

// Look-up table parameters
//

`define DSP58_ADDR_N  50
`define DSP58_ADDR_SZ 32
`define DSP58_DATA_SZ 120

// Attribute addresses
//

`define DSP58__ACASCREG    32'h00000000
`define DSP58__ACASCREG_SZ 32

`define DSP58__ADREG    32'h00000001
`define DSP58__ADREG_SZ 32

`define DSP58__ALUMODEREG    32'h00000002
`define DSP58__ALUMODEREG_SZ 32

`define DSP58__AMULTSEL    32'h00000003
`define DSP58__AMULTSEL_SZ 16

`define DSP58__AREG    32'h00000004
`define DSP58__AREG_SZ 32

`define DSP58__AUTORESET_PATDET    32'h00000005
`define DSP58__AUTORESET_PATDET_SZ 120

`define DSP58__AUTORESET_PRIORITY    32'h00000006
`define DSP58__AUTORESET_PRIORITY_SZ 40

`define DSP58__A_INPUT    32'h00000007
`define DSP58__A_INPUT_SZ 56

`define DSP58__BCASCREG    32'h00000008
`define DSP58__BCASCREG_SZ 32

`define DSP58__BMULTSEL    32'h00000009
`define DSP58__BMULTSEL_SZ 16

`define DSP58__BREG    32'h0000000a
`define DSP58__BREG_SZ 32

`define DSP58__B_INPUT    32'h0000000b
`define DSP58__B_INPUT_SZ 56

`define DSP58__CARRYINREG    32'h0000000c
`define DSP58__CARRYINREG_SZ 32

`define DSP58__CARRYINSELREG    32'h0000000d
`define DSP58__CARRYINSELREG_SZ 32

`define DSP58__CREG    32'h0000000e
`define DSP58__CREG_SZ 32

`define DSP58__DREG    32'h0000000f
`define DSP58__DREG_SZ 32

`define DSP58__DSP_MODE    32'h00000010
`define DSP58__DSP_MODE_SZ 40

`define DSP58__INMODEREG    32'h00000011
`define DSP58__INMODEREG_SZ 32

`define DSP58__IS_ALUMODE_INVERTED    32'h00000012
`define DSP58__IS_ALUMODE_INVERTED_SZ 4

`define DSP58__IS_ASYNC_RST_INVERTED    32'h00000013
`define DSP58__IS_ASYNC_RST_INVERTED_SZ 1

`define DSP58__IS_CARRYIN_INVERTED    32'h00000014
`define DSP58__IS_CARRYIN_INVERTED_SZ 1

`define DSP58__IS_CLK_INVERTED    32'h00000015
`define DSP58__IS_CLK_INVERTED_SZ 1

`define DSP58__IS_INMODE_INVERTED    32'h00000016
`define DSP58__IS_INMODE_INVERTED_SZ 5

`define DSP58__IS_NEGATE_INVERTED    32'h00000017
`define DSP58__IS_NEGATE_INVERTED_SZ 3

`define DSP58__IS_OPMODE_INVERTED    32'h00000018
`define DSP58__IS_OPMODE_INVERTED_SZ 9

`define DSP58__IS_RSTALLCARRYIN_INVERTED    32'h00000019
`define DSP58__IS_RSTALLCARRYIN_INVERTED_SZ 1

`define DSP58__IS_RSTALUMODE_INVERTED    32'h0000001a
`define DSP58__IS_RSTALUMODE_INVERTED_SZ 1

`define DSP58__IS_RSTA_INVERTED    32'h0000001b
`define DSP58__IS_RSTA_INVERTED_SZ 1

`define DSP58__IS_RSTB_INVERTED    32'h0000001c
`define DSP58__IS_RSTB_INVERTED_SZ 1

`define DSP58__IS_RSTCTRL_INVERTED    32'h0000001d
`define DSP58__IS_RSTCTRL_INVERTED_SZ 1

`define DSP58__IS_RSTC_INVERTED    32'h0000001e
`define DSP58__IS_RSTC_INVERTED_SZ 1

`define DSP58__IS_RSTD_INVERTED    32'h0000001f
`define DSP58__IS_RSTD_INVERTED_SZ 1

`define DSP58__IS_RSTINMODE_INVERTED    32'h00000020
`define DSP58__IS_RSTINMODE_INVERTED_SZ 1

`define DSP58__IS_RSTM_INVERTED    32'h00000021
`define DSP58__IS_RSTM_INVERTED_SZ 1

`define DSP58__IS_RSTP_INVERTED    32'h00000022
`define DSP58__IS_RSTP_INVERTED_SZ 1

`define DSP58__MASK    32'h00000023
`define DSP58__MASK_SZ 58

`define DSP58__MREG    32'h00000024
`define DSP58__MREG_SZ 32

`define DSP58__OPMODEREG    32'h00000025
`define DSP58__OPMODEREG_SZ 32

`define DSP58__PATTERN    32'h00000026
`define DSP58__PATTERN_SZ 58

`define DSP58__PREADDINSEL    32'h00000027
`define DSP58__PREADDINSEL_SZ 8

`define DSP58__PREG    32'h00000028
`define DSP58__PREG_SZ 32

`define DSP58__RESET_MODE    32'h00000029
`define DSP58__RESET_MODE_SZ 40

`define DSP58__RND    32'h0000002a
`define DSP58__RND_SZ 58

`define DSP58__SEL_MASK    32'h0000002b
`define DSP58__SEL_MASK_SZ 112

`define DSP58__SEL_PATTERN    32'h0000002c
`define DSP58__SEL_PATTERN_SZ 56

`define DSP58__USE_MULT    32'h0000002d
`define DSP58__USE_MULT_SZ 64

`define DSP58__USE_PATTERN_DETECT    32'h0000002e
`define DSP58__USE_PATTERN_DETECT_SZ 72

`define DSP58__USE_SIMD    32'h0000002f
`define DSP58__USE_SIMD_SZ 48

`define DSP58__USE_WIDEXOR    32'h00000030
`define DSP58__USE_WIDEXOR_SZ 40

`define DSP58__XORSIMD    32'h00000031
`define DSP58__XORSIMD_SZ 120

`endif  // B_DSP58_DEFINES_VH