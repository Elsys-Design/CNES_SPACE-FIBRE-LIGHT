`include "B_DSP_FP_OUTPUT_defines.vh"

reg [`DSP_FP_OUTPUT_DATA_SZ-1:0] ATTR [0:`DSP_FP_OUTPUT_ADDR_N-1];
reg [`DSP_FP_OUTPUT__FPA_PREG_SZ-1:0] FPA_PREG_REG = FPA_PREG;
reg [`DSP_FP_OUTPUT__FPM_PREG_SZ-1:0] FPM_PREG_REG = FPM_PREG;
reg IS_RSTFPA_INVERTED_REG = IS_RSTFPA_INVERTED;
reg IS_RSTFPM_INVERTED_REG = IS_RSTFPM_INVERTED;
reg [`DSP_FP_OUTPUT__PCOUTSEL_SZ:1] PCOUTSEL_REG = PCOUTSEL;
reg [`DSP_FP_OUTPUT__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;
reg [`DSP_FP_OUTPUT__USE_MULT_SZ:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_FP_OUTPUT__FPA_PREG] = FPA_PREG;
  ATTR[`DSP_FP_OUTPUT__FPM_PREG] = FPM_PREG;
  ATTR[`DSP_FP_OUTPUT__IS_RSTFPA_INVERTED] = IS_RSTFPA_INVERTED;
  ATTR[`DSP_FP_OUTPUT__IS_RSTFPM_INVERTED] = IS_RSTFPM_INVERTED;
  ATTR[`DSP_FP_OUTPUT__PCOUTSEL] = PCOUTSEL;
  ATTR[`DSP_FP_OUTPUT__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_FP_OUTPUT__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  FPA_PREG_REG = ATTR[`DSP_FP_OUTPUT__FPA_PREG];
  FPM_PREG_REG = ATTR[`DSP_FP_OUTPUT__FPM_PREG];
  IS_RSTFPA_INVERTED_REG = ATTR[`DSP_FP_OUTPUT__IS_RSTFPA_INVERTED];
  IS_RSTFPM_INVERTED_REG = ATTR[`DSP_FP_OUTPUT__IS_RSTFPM_INVERTED];
  PCOUTSEL_REG = ATTR[`DSP_FP_OUTPUT__PCOUTSEL];
  RESET_MODE_REG = ATTR[`DSP_FP_OUTPUT__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_FP_OUTPUT__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FP_OUTPUT_ADDR_SZ-1:0] addr;
  input  [`DSP_FP_OUTPUT_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FP_OUTPUT_DATA_SZ-1:0] read_attr;
  input  [`DSP_FP_OUTPUT_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
