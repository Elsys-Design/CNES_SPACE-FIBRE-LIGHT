// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_BUFGCTRL_DEFINES_VH
`else
`define B_BUFGCTRL_DEFINES_VH

// Look-up table parameters
//

`define BUFGCTRL_ADDR_N  15
`define BUFGCTRL_ADDR_SZ 32
`define BUFGCTRL_DATA_SZ 144

// Attribute addresses
//

`define BUFGCTRL__CE_TYPE_CE0    32'h00000000
`define BUFGCTRL__CE_TYPE_CE0_SZ 64

`define BUFGCTRL__CE_TYPE_CE1    32'h00000001
`define BUFGCTRL__CE_TYPE_CE1_SZ 64

`define BUFGCTRL__INIT_OUT    32'h00000002
`define BUFGCTRL__INIT_OUT_SZ 32

`define BUFGCTRL__IS_CE0_INVERTED    32'h00000003
`define BUFGCTRL__IS_CE0_INVERTED_SZ 1

`define BUFGCTRL__IS_CE1_INVERTED    32'h00000004
`define BUFGCTRL__IS_CE1_INVERTED_SZ 1

`define BUFGCTRL__IS_I0_INVERTED    32'h00000005
`define BUFGCTRL__IS_I0_INVERTED_SZ 1

`define BUFGCTRL__IS_I1_INVERTED    32'h00000006
`define BUFGCTRL__IS_I1_INVERTED_SZ 1

`define BUFGCTRL__IS_IGNORE0_INVERTED    32'h00000007
`define BUFGCTRL__IS_IGNORE0_INVERTED_SZ 1

`define BUFGCTRL__IS_IGNORE1_INVERTED    32'h00000008
`define BUFGCTRL__IS_IGNORE1_INVERTED_SZ 1

`define BUFGCTRL__IS_S0_INVERTED    32'h00000009
`define BUFGCTRL__IS_S0_INVERTED_SZ 1

`define BUFGCTRL__IS_S1_INVERTED    32'h0000000a
`define BUFGCTRL__IS_S1_INVERTED_SZ 1

`define BUFGCTRL__PRESELECT_I0    32'h0000000b
`define BUFGCTRL__PRESELECT_I0_SZ 40

`define BUFGCTRL__PRESELECT_I1    32'h0000000c
`define BUFGCTRL__PRESELECT_I1_SZ 40

`define BUFGCTRL__SIM_DEVICE    32'h0000000d
`define BUFGCTRL__SIM_DEVICE_SZ 144

`define BUFGCTRL__STARTUP_SYNC    32'h0000000e
`define BUFGCTRL__STARTUP_SYNC_SZ 40

`endif  // B_BUFGCTRL_DEFINES_VH
