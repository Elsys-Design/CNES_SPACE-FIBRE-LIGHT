`include "B_MBUFGCE_DIV_defines.vh"

reg [`MBUFGCE_DIV_DATA_SZ-1:0] ATTR [0:`MBUFGCE_DIV_ADDR_N-1];
reg [`MBUFGCE_DIV__BUFGCE_DIVIDE_SZ-1:0] BUFGCE_DIVIDE_REG = BUFGCE_DIVIDE;
reg [`MBUFGCE_DIV__CE_TYPE_SZ:1] CE_TYPE_REG = CE_TYPE;
reg [`MBUFGCE_DIV__HARDSYNC_CLR_SZ:1] HARDSYNC_CLR_REG = HARDSYNC_CLR;
reg IS_CE_INVERTED_REG = IS_CE_INVERTED;
reg IS_CLR_INVERTED_REG = IS_CLR_INVERTED;
reg IS_I_INVERTED_REG = IS_I_INVERTED;
reg [`MBUFGCE_DIV__MODE_SZ:1] MODE_REG = MODE;
reg [`MBUFGCE_DIV__STARTUP_SYNC_SZ:1] STARTUP_SYNC_REG = STARTUP_SYNC;

initial begin
  ATTR[`MBUFGCE_DIV__BUFGCE_DIVIDE] = BUFGCE_DIVIDE;
  ATTR[`MBUFGCE_DIV__CE_TYPE] = CE_TYPE;
  ATTR[`MBUFGCE_DIV__HARDSYNC_CLR] = HARDSYNC_CLR;
  ATTR[`MBUFGCE_DIV__IS_CE_INVERTED] = IS_CE_INVERTED;
  ATTR[`MBUFGCE_DIV__IS_CLR_INVERTED] = IS_CLR_INVERTED;
  ATTR[`MBUFGCE_DIV__IS_I_INVERTED] = IS_I_INVERTED;
  ATTR[`MBUFGCE_DIV__MODE] = MODE;
  ATTR[`MBUFGCE_DIV__STARTUP_SYNC] = STARTUP_SYNC;
end

always @(trig_attr) begin
  BUFGCE_DIVIDE_REG = ATTR[`MBUFGCE_DIV__BUFGCE_DIVIDE];
  CE_TYPE_REG = ATTR[`MBUFGCE_DIV__CE_TYPE];
  HARDSYNC_CLR_REG = ATTR[`MBUFGCE_DIV__HARDSYNC_CLR];
  IS_CE_INVERTED_REG = ATTR[`MBUFGCE_DIV__IS_CE_INVERTED];
  IS_CLR_INVERTED_REG = ATTR[`MBUFGCE_DIV__IS_CLR_INVERTED];
  IS_I_INVERTED_REG = ATTR[`MBUFGCE_DIV__IS_I_INVERTED];
  MODE_REG = ATTR[`MBUFGCE_DIV__MODE];
  STARTUP_SYNC_REG = ATTR[`MBUFGCE_DIV__STARTUP_SYNC];
end

// procedures to override, read attribute values

task write_attr;
  input  [`MBUFGCE_DIV_ADDR_SZ-1:0] addr;
  input  [`MBUFGCE_DIV_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`MBUFGCE_DIV_DATA_SZ-1:0] read_attr;
  input  [`MBUFGCE_DIV_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
