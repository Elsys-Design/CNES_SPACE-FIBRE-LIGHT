// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_FP_INREG_DEFINES_VH
`else
`define B_DSP_FP_INREG_DEFINES_VH

// Look-up table parameters
//

`define DSP_FP_INREG_ADDR_N  12
`define DSP_FP_INREG_ADDR_SZ 32
`define DSP_FP_INREG_DATA_SZ 56

// Attribute addresses
//

`define DSP_FP_INREG__ACASCREG    32'h00000000
`define DSP_FP_INREG__ACASCREG_SZ 32

`define DSP_FP_INREG__AREG    32'h00000001
`define DSP_FP_INREG__AREG_SZ 32

`define DSP_FP_INREG__A_FPTYPE    32'h00000002
`define DSP_FP_INREG__A_FPTYPE_SZ 24

`define DSP_FP_INREG__A_INPUT    32'h00000003
`define DSP_FP_INREG__A_INPUT_SZ 56

`define DSP_FP_INREG__BCASCSEL    32'h00000004
`define DSP_FP_INREG__BCASCSEL_SZ 8

`define DSP_FP_INREG__B_D_FPTYPE    32'h00000005
`define DSP_FP_INREG__B_D_FPTYPE_SZ 24

`define DSP_FP_INREG__B_INPUT    32'h00000006
`define DSP_FP_INREG__B_INPUT_SZ 56

`define DSP_FP_INREG__FPBREG    32'h00000007
`define DSP_FP_INREG__FPBREG_SZ 32

`define DSP_FP_INREG__FPDREG    32'h00000008
`define DSP_FP_INREG__FPDREG_SZ 32

`define DSP_FP_INREG__IS_RSTA_INVERTED    32'h00000009
`define DSP_FP_INREG__IS_RSTA_INVERTED_SZ 1

`define DSP_FP_INREG__IS_RSTB_INVERTED    32'h0000000a
`define DSP_FP_INREG__IS_RSTB_INVERTED_SZ 1

`define DSP_FP_INREG__RESET_MODE    32'h0000000b
`define DSP_FP_INREG__RESET_MODE_SZ 40

`endif  // B_DSP_FP_INREG_DEFINES_VH