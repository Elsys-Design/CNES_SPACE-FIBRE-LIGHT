// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_MMCME5_DEFINES_VH
`else
`define B_MMCME5_DEFINES_VH

// Look-up table parameters
//

`define MMCME5_ADDR_N  67
`define MMCME5_ADDR_SZ 32
`define MMCME5_DATA_SZ 88

// Attribute addresses
//

`define MMCME5__BANDWIDTH    32'h00000000
`define MMCME5__BANDWIDTH_SZ 72

`define MMCME5__CLKFBOUT_FRACT    32'h00000001
`define MMCME5__CLKFBOUT_FRACT_SZ 32

`define MMCME5__CLKFBOUT_MULT    32'h00000002
`define MMCME5__CLKFBOUT_MULT_SZ 32

`define MMCME5__CLKFBOUT_PHASE    32'h00000003
`define MMCME5__CLKFBOUT_PHASE_SZ 64

`define MMCME5__CLKIN1_PERIOD    32'h00000004
`define MMCME5__CLKIN1_PERIOD_SZ 64

`define MMCME5__CLKIN2_PERIOD    32'h00000005
`define MMCME5__CLKIN2_PERIOD_SZ 64

`define MMCME5__CLKIN_FREQ_MAX    32'h00000006
`define MMCME5__CLKIN_FREQ_MAX_SZ 64

`define MMCME5__CLKIN_FREQ_MIN    32'h00000007
`define MMCME5__CLKIN_FREQ_MIN_SZ 64

`define MMCME5__CLKOUT0_DIVIDE    32'h00000008
`define MMCME5__CLKOUT0_DIVIDE_SZ 32

`define MMCME5__CLKOUT0_DUTY_CYCLE    32'h00000009
`define MMCME5__CLKOUT0_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT0_PHASE    32'h0000000a
`define MMCME5__CLKOUT0_PHASE_SZ 64

`define MMCME5__CLKOUT0_PHASE_CTRL    32'h0000000b
`define MMCME5__CLKOUT0_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT1_DIVIDE    32'h0000000c
`define MMCME5__CLKOUT1_DIVIDE_SZ 32

`define MMCME5__CLKOUT1_DUTY_CYCLE    32'h0000000d
`define MMCME5__CLKOUT1_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT1_PHASE    32'h0000000e
`define MMCME5__CLKOUT1_PHASE_SZ 64

`define MMCME5__CLKOUT1_PHASE_CTRL    32'h0000000f
`define MMCME5__CLKOUT1_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT2_DIVIDE    32'h00000010
`define MMCME5__CLKOUT2_DIVIDE_SZ 32

`define MMCME5__CLKOUT2_DUTY_CYCLE    32'h00000011
`define MMCME5__CLKOUT2_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT2_PHASE    32'h00000012
`define MMCME5__CLKOUT2_PHASE_SZ 64

`define MMCME5__CLKOUT2_PHASE_CTRL    32'h00000013
`define MMCME5__CLKOUT2_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT3_DIVIDE    32'h00000014
`define MMCME5__CLKOUT3_DIVIDE_SZ 32

`define MMCME5__CLKOUT3_DUTY_CYCLE    32'h00000015
`define MMCME5__CLKOUT3_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT3_PHASE    32'h00000016
`define MMCME5__CLKOUT3_PHASE_SZ 64

`define MMCME5__CLKOUT3_PHASE_CTRL    32'h00000017
`define MMCME5__CLKOUT3_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT4_DIVIDE    32'h00000018
`define MMCME5__CLKOUT4_DIVIDE_SZ 32

`define MMCME5__CLKOUT4_DUTY_CYCLE    32'h00000019
`define MMCME5__CLKOUT4_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT4_PHASE    32'h0000001a
`define MMCME5__CLKOUT4_PHASE_SZ 64

`define MMCME5__CLKOUT4_PHASE_CTRL    32'h0000001b
`define MMCME5__CLKOUT4_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT5_DIVIDE    32'h0000001c
`define MMCME5__CLKOUT5_DIVIDE_SZ 32

`define MMCME5__CLKOUT5_DUTY_CYCLE    32'h0000001d
`define MMCME5__CLKOUT5_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT5_PHASE    32'h0000001e
`define MMCME5__CLKOUT5_PHASE_SZ 64

`define MMCME5__CLKOUT5_PHASE_CTRL    32'h0000001f
`define MMCME5__CLKOUT5_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUT6_DIVIDE    32'h00000020
`define MMCME5__CLKOUT6_DIVIDE_SZ 32

`define MMCME5__CLKOUT6_DUTY_CYCLE    32'h00000021
`define MMCME5__CLKOUT6_DUTY_CYCLE_SZ 64

`define MMCME5__CLKOUT6_PHASE    32'h00000022
`define MMCME5__CLKOUT6_PHASE_SZ 64

`define MMCME5__CLKOUT6_PHASE_CTRL    32'h00000023
`define MMCME5__CLKOUT6_PHASE_CTRL_SZ 2

`define MMCME5__CLKOUTFB_PHASE_CTRL    32'h00000024
`define MMCME5__CLKOUTFB_PHASE_CTRL_SZ 2

`define MMCME5__CLKPFD_FREQ_MAX    32'h00000025
`define MMCME5__CLKPFD_FREQ_MAX_SZ 64

`define MMCME5__CLKPFD_FREQ_MIN    32'h00000026
`define MMCME5__CLKPFD_FREQ_MIN_SZ 64

`define MMCME5__COMPENSATION    32'h00000027
`define MMCME5__COMPENSATION_SZ 64

`define MMCME5__DESKEW_DELAY1    32'h00000028
`define MMCME5__DESKEW_DELAY1_SZ 32

`define MMCME5__DESKEW_DELAY2    32'h00000029
`define MMCME5__DESKEW_DELAY2_SZ 32

`define MMCME5__DESKEW_DELAY_EN1    32'h0000002a
`define MMCME5__DESKEW_DELAY_EN1_SZ 40

`define MMCME5__DESKEW_DELAY_EN2    32'h0000002b
`define MMCME5__DESKEW_DELAY_EN2_SZ 40

`define MMCME5__DESKEW_DELAY_PATH1    32'h0000002c
`define MMCME5__DESKEW_DELAY_PATH1_SZ 40

`define MMCME5__DESKEW_DELAY_PATH2    32'h0000002d
`define MMCME5__DESKEW_DELAY_PATH2_SZ 40

`define MMCME5__DIVCLK_DIVIDE    32'h0000002e
`define MMCME5__DIVCLK_DIVIDE_SZ 32

`define MMCME5__IS_CLKFB1_DESKEW_INVERTED    32'h0000002f
`define MMCME5__IS_CLKFB1_DESKEW_INVERTED_SZ 1

`define MMCME5__IS_CLKFB2_DESKEW_INVERTED    32'h00000030
`define MMCME5__IS_CLKFB2_DESKEW_INVERTED_SZ 1

`define MMCME5__IS_CLKFBIN_INVERTED    32'h00000031
`define MMCME5__IS_CLKFBIN_INVERTED_SZ 1

`define MMCME5__IS_CLKIN1_DESKEW_INVERTED    32'h00000032
`define MMCME5__IS_CLKIN1_DESKEW_INVERTED_SZ 1

`define MMCME5__IS_CLKIN1_INVERTED    32'h00000033
`define MMCME5__IS_CLKIN1_INVERTED_SZ 1

`define MMCME5__IS_CLKIN2_DESKEW_INVERTED    32'h00000034
`define MMCME5__IS_CLKIN2_DESKEW_INVERTED_SZ 1

`define MMCME5__IS_CLKIN2_INVERTED    32'h00000035
`define MMCME5__IS_CLKIN2_INVERTED_SZ 1

`define MMCME5__IS_CLKINSEL_INVERTED    32'h00000036
`define MMCME5__IS_CLKINSEL_INVERTED_SZ 1

`define MMCME5__IS_PSEN_INVERTED    32'h00000037
`define MMCME5__IS_PSEN_INVERTED_SZ 1

`define MMCME5__IS_PSINCDEC_INVERTED    32'h00000038
`define MMCME5__IS_PSINCDEC_INVERTED_SZ 1

`define MMCME5__IS_PWRDWN_INVERTED    32'h00000039
`define MMCME5__IS_PWRDWN_INVERTED_SZ 1

`define MMCME5__IS_RST_INVERTED    32'h0000003a
`define MMCME5__IS_RST_INVERTED_SZ 1

`define MMCME5__LOCK_WAIT    32'h0000003b
`define MMCME5__LOCK_WAIT_SZ 40

`define MMCME5__REF_JITTER1    32'h0000003c
`define MMCME5__REF_JITTER1_SZ 64

`define MMCME5__REF_JITTER2    32'h0000003d
`define MMCME5__REF_JITTER2_SZ 64

`define MMCME5__SS_EN    32'h0000003e
`define MMCME5__SS_EN_SZ 40

`define MMCME5__SS_MODE    32'h0000003f
`define MMCME5__SS_MODE_SZ 88

`define MMCME5__SS_MOD_PERIOD    32'h00000040
`define MMCME5__SS_MOD_PERIOD_SZ 32

`define MMCME5__VCOCLK_FREQ_MAX    32'h00000041
`define MMCME5__VCOCLK_FREQ_MAX_SZ 64

`define MMCME5__VCOCLK_FREQ_MIN    32'h00000042
`define MMCME5__VCOCLK_FREQ_MIN_SZ 64

`endif  // B_MMCME5_DEFINES_VH