-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 18/07/2025
--
-- Description : This module implements the parallel loopback function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_parallel_loopback is
    port (
      CLK                      : in  std_logic;                                   --! Clock generated by HSSL IP
      RST_N                    : in  std_logic;                                   --! Global reset. Active low
      -- ppl_64_lane_ctrl_word_insert (PLCWI) interface
      DATA_TX_PLCWI            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CARAC_PLCWI      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLCWI           : in  std_logic;                                   --! Data ready flag
      -- ppl_64_rx_sync_fsm (PLRSF) interface
      DATA_TX_PLRSF            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CARAC_PLRSF      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLRSF           : in  std_logic;                                   --! Data ready flag
      LOSS_OF_SIGNAL_PLRSF     : in  std_logic;                                   --! Loss of signal flag from PLRSF
      -- ppl_64_skip_insertion (PLSI) interface
      WAIT_SEND_DATA_PLSI      : in  std_logic;                                   --! Wait send data signal for SKIP insertion
      -- ppl_64_lane_ctrl_word_detection (PLCWD) interface
      DATA_RX_PLPL             : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit Data
      VALID_K_CHARAC_PLPL      : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit Valid K character
      DATA_RDY_PLPL            : out std_logic;                                   --! Data ready flag
      LOSS_OF_SIGNAL_PLPL      : out std_logic;                                   --! Loss of signal flag from PLPL 
      -- MIB interface
      PARALLEL_LOOPBACK_EN_MIB : in  std_logic                                    --! Enable or disable the parallel loopback
    );
end ppl_64_parallel_loopback;

architecture rtl of ppl_64_parallel_loopback is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
signal wait_send_data_r                : std_logic;
signal wait_send_data_rr               : std_logic;
signal wait_send_data_rrr              : std_logic;

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_delay_wait_send_data
  --! Delays the wait_send_data signal
  ---------------------------------------------------------
  p_delay_wait_send_data : process(CLK, RST_N)
  begin
    if RST_N = '0' then
      wait_send_data_r   <= '0';
      wait_send_data_rr  <= '0';
      wait_send_data_rrr <= '0';
    elsif rising_edge(CLK) then
      wait_send_data_r   <= WAIT_SEND_DATA_PLSI;
      wait_send_data_rr  <= wait_send_data_r;
      wait_send_data_rrr <= wait_send_data_rr;
    end if;
  end process p_delay_wait_send_data;

  -- Allows a parallel loopback into the LANE layer
  DATA_RX_PLPL        <= DATA_TX_PLCWI                                    when PARALLEL_LOOPBACK_EN_MIB = '1' else DATA_TX_PLRSF;
  VALID_K_CHARAC_PLPL <= VALID_K_CARAC_PLCWI                              when PARALLEL_LOOPBACK_EN_MIB = '1' else VALID_K_CARAC_PLRSF;
  DATA_RDY_PLPL       <= (DATA_RDY_PLCWI and not(wait_send_data_rrr) )    when PARALLEL_LOOPBACK_EN_MIB = '1' else DATA_RDY_PLRSF;
  LOSS_OF_SIGNAL_PLPL <= '0'                                              when PARALLEL_LOOPBACK_EN_MIB = '1' else LOSS_OF_SIGNAL_PLRSF;
end architecture rtl;
