// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_ILKNE4_DEFINES_VH
`else
`define B_ILKNE4_DEFINES_VH

// Look-up table parameters
//

`define ILKNE4_ADDR_N  26
`define ILKNE4_ADDR_SZ 32
`define ILKNE4_DATA_SZ 152

// Attribute addresses
//

`define ILKNE4__BYPASS    32'h00000000
`define ILKNE4__BYPASS_SZ 40

`define ILKNE4__CTL_RX_BURSTMAX    32'h00000001
`define ILKNE4__CTL_RX_BURSTMAX_SZ 2

`define ILKNE4__CTL_RX_CHAN_EXT    32'h00000002
`define ILKNE4__CTL_RX_CHAN_EXT_SZ 2

`define ILKNE4__CTL_RX_LAST_LANE    32'h00000003
`define ILKNE4__CTL_RX_LAST_LANE_SZ 4

`define ILKNE4__CTL_RX_MFRAMELEN_MINUS1    32'h00000004
`define ILKNE4__CTL_RX_MFRAMELEN_MINUS1_SZ 16

`define ILKNE4__CTL_RX_PACKET_MODE    32'h00000005
`define ILKNE4__CTL_RX_PACKET_MODE_SZ 40

`define ILKNE4__CTL_RX_RETRANS_MULT    32'h00000006
`define ILKNE4__CTL_RX_RETRANS_MULT_SZ 3

`define ILKNE4__CTL_RX_RETRANS_RETRY    32'h00000007
`define ILKNE4__CTL_RX_RETRANS_RETRY_SZ 4

`define ILKNE4__CTL_RX_RETRANS_TIMER1    32'h00000008
`define ILKNE4__CTL_RX_RETRANS_TIMER1_SZ 16

`define ILKNE4__CTL_RX_RETRANS_TIMER2    32'h00000009
`define ILKNE4__CTL_RX_RETRANS_TIMER2_SZ 16

`define ILKNE4__CTL_RX_RETRANS_WDOG    32'h0000000a
`define ILKNE4__CTL_RX_RETRANS_WDOG_SZ 12

`define ILKNE4__CTL_RX_RETRANS_WRAP_TIMER    32'h0000000b
`define ILKNE4__CTL_RX_RETRANS_WRAP_TIMER_SZ 8

`define ILKNE4__CTL_TEST_MODE_PIN_CHAR    32'h0000000c
`define ILKNE4__CTL_TEST_MODE_PIN_CHAR_SZ 40

`define ILKNE4__CTL_TX_BURSTMAX    32'h0000000d
`define ILKNE4__CTL_TX_BURSTMAX_SZ 2

`define ILKNE4__CTL_TX_BURSTSHORT    32'h0000000e
`define ILKNE4__CTL_TX_BURSTSHORT_SZ 3

`define ILKNE4__CTL_TX_CHAN_EXT    32'h0000000f
`define ILKNE4__CTL_TX_CHAN_EXT_SZ 2

`define ILKNE4__CTL_TX_DISABLE_SKIPWORD    32'h00000010
`define ILKNE4__CTL_TX_DISABLE_SKIPWORD_SZ 40

`define ILKNE4__CTL_TX_FC_CALLEN    32'h00000011
`define ILKNE4__CTL_TX_FC_CALLEN_SZ 4

`define ILKNE4__CTL_TX_LAST_LANE    32'h00000012
`define ILKNE4__CTL_TX_LAST_LANE_SZ 4

`define ILKNE4__CTL_TX_MFRAMELEN_MINUS1    32'h00000013
`define ILKNE4__CTL_TX_MFRAMELEN_MINUS1_SZ 16

`define ILKNE4__CTL_TX_RETRANS_DEPTH    32'h00000014
`define ILKNE4__CTL_TX_RETRANS_DEPTH_SZ 14

`define ILKNE4__CTL_TX_RETRANS_MULT    32'h00000015
`define ILKNE4__CTL_TX_RETRANS_MULT_SZ 3

`define ILKNE4__CTL_TX_RETRANS_RAM_BANKS    32'h00000016
`define ILKNE4__CTL_TX_RETRANS_RAM_BANKS_SZ 2

`define ILKNE4__MODE    32'h00000017
`define ILKNE4__MODE_SZ 40

`define ILKNE4__SIM_DEVICE    32'h00000018
`define ILKNE4__SIM_DEVICE_SZ 152

`define ILKNE4__TEST_MODE_PIN_CHAR    32'h00000019
`define ILKNE4__TEST_MODE_PIN_CHAR_SZ 40

`endif  // B_ILKNE4_DEFINES_VH