`include "B_DSP_A_B_DATA58_defines.vh"

reg [`DSP_A_B_DATA58_DATA_SZ-1:0] ATTR [0:`DSP_A_B_DATA58_ADDR_N-1];
reg [`DSP_A_B_DATA58__ACASCREG_SZ-1:0] ACASCREG_REG = ACASCREG;
reg [`DSP_A_B_DATA58__AMULTSEL_SZ:1] AMULTSEL_REG = AMULTSEL;
reg [`DSP_A_B_DATA58__AREG_SZ-1:0] AREG_REG = AREG;
reg [`DSP_A_B_DATA58__A_INPUT_SZ:1] A_INPUT_REG = A_INPUT;
reg [`DSP_A_B_DATA58__BCASCREG_SZ-1:0] BCASCREG_REG = BCASCREG;
reg [`DSP_A_B_DATA58__BMULTSEL_SZ:1] BMULTSEL_REG = BMULTSEL;
reg [`DSP_A_B_DATA58__BREG_SZ-1:0] BREG_REG = BREG;
reg [`DSP_A_B_DATA58__B_INPUT_SZ:1] B_INPUT_REG = B_INPUT;
reg [`DSP_A_B_DATA58__DSP_MODE_SZ:1] DSP_MODE_REG = DSP_MODE;
reg IS_RSTA_INVERTED_REG = IS_RSTA_INVERTED;
reg IS_RSTB_INVERTED_REG = IS_RSTB_INVERTED;
reg [`DSP_A_B_DATA58__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;

initial begin
  ATTR[`DSP_A_B_DATA58__ACASCREG] = ACASCREG;
  ATTR[`DSP_A_B_DATA58__AMULTSEL] = AMULTSEL;
  ATTR[`DSP_A_B_DATA58__AREG] = AREG;
  ATTR[`DSP_A_B_DATA58__A_INPUT] = A_INPUT;
  ATTR[`DSP_A_B_DATA58__BCASCREG] = BCASCREG;
  ATTR[`DSP_A_B_DATA58__BMULTSEL] = BMULTSEL;
  ATTR[`DSP_A_B_DATA58__BREG] = BREG;
  ATTR[`DSP_A_B_DATA58__B_INPUT] = B_INPUT;
  ATTR[`DSP_A_B_DATA58__DSP_MODE] = DSP_MODE;
  ATTR[`DSP_A_B_DATA58__IS_RSTA_INVERTED] = IS_RSTA_INVERTED;
  ATTR[`DSP_A_B_DATA58__IS_RSTB_INVERTED] = IS_RSTB_INVERTED;
  ATTR[`DSP_A_B_DATA58__RESET_MODE] = RESET_MODE;
end

always @(*) begin
  ACASCREG_REG = ATTR[`DSP_A_B_DATA58__ACASCREG];
  AMULTSEL_REG = ATTR[`DSP_A_B_DATA58__AMULTSEL];
  AREG_REG = ATTR[`DSP_A_B_DATA58__AREG];
  A_INPUT_REG = ATTR[`DSP_A_B_DATA58__A_INPUT];
  BCASCREG_REG = ATTR[`DSP_A_B_DATA58__BCASCREG];
  BMULTSEL_REG = ATTR[`DSP_A_B_DATA58__BMULTSEL];
  BREG_REG = ATTR[`DSP_A_B_DATA58__BREG];
  B_INPUT_REG = ATTR[`DSP_A_B_DATA58__B_INPUT];
  DSP_MODE_REG = ATTR[`DSP_A_B_DATA58__DSP_MODE];
  IS_RSTA_INVERTED_REG = ATTR[`DSP_A_B_DATA58__IS_RSTA_INVERTED];
  IS_RSTB_INVERTED_REG = ATTR[`DSP_A_B_DATA58__IS_RSTB_INVERTED];
  RESET_MODE_REG = ATTR[`DSP_A_B_DATA58__RESET_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_A_B_DATA58_ADDR_SZ-1:0] addr;
  input  [`DSP_A_B_DATA58_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_A_B_DATA58_DATA_SZ-1:0] read_attr;
  input  [`DSP_A_B_DATA58_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
