// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_PLLE4_BASE_DEFINES_VH
`else
`define B_PLLE4_BASE_DEFINES_VH

// Look-up table parameters
//

`define PLLE4_BASE_ADDR_N  17
`define PLLE4_BASE_ADDR_SZ 32
`define PLLE4_BASE_DATA_SZ 64

// Attribute addresses
//

`define PLLE4_BASE__CLKFBOUT_MULT    32'h00000000
`define PLLE4_BASE__CLKFBOUT_MULT_SZ 32

`define PLLE4_BASE__CLKFBOUT_PHASE    32'h00000001
`define PLLE4_BASE__CLKFBOUT_PHASE_SZ 64

`define PLLE4_BASE__CLKIN_PERIOD    32'h00000002
`define PLLE4_BASE__CLKIN_PERIOD_SZ 64

`define PLLE4_BASE__CLKOUT0_DIVIDE    32'h00000003
`define PLLE4_BASE__CLKOUT0_DIVIDE_SZ 32

`define PLLE4_BASE__CLKOUT0_DUTY_CYCLE    32'h00000004
`define PLLE4_BASE__CLKOUT0_DUTY_CYCLE_SZ 64

`define PLLE4_BASE__CLKOUT0_PHASE    32'h00000005
`define PLLE4_BASE__CLKOUT0_PHASE_SZ 64

`define PLLE4_BASE__CLKOUT1_DIVIDE    32'h00000006
`define PLLE4_BASE__CLKOUT1_DIVIDE_SZ 32

`define PLLE4_BASE__CLKOUT1_DUTY_CYCLE    32'h00000007
`define PLLE4_BASE__CLKOUT1_DUTY_CYCLE_SZ 64

`define PLLE4_BASE__CLKOUT1_PHASE    32'h00000008
`define PLLE4_BASE__CLKOUT1_PHASE_SZ 64

`define PLLE4_BASE__CLKOUTPHY_MODE    32'h00000009
`define PLLE4_BASE__CLKOUTPHY_MODE_SZ 64

`define PLLE4_BASE__DIVCLK_DIVIDE    32'h0000000a
`define PLLE4_BASE__DIVCLK_DIVIDE_SZ 32

`define PLLE4_BASE__IS_CLKFBIN_INVERTED    32'h0000000b
`define PLLE4_BASE__IS_CLKFBIN_INVERTED_SZ 1

`define PLLE4_BASE__IS_CLKIN_INVERTED    32'h0000000c
`define PLLE4_BASE__IS_CLKIN_INVERTED_SZ 1

`define PLLE4_BASE__IS_PWRDWN_INVERTED    32'h0000000d
`define PLLE4_BASE__IS_PWRDWN_INVERTED_SZ 1

`define PLLE4_BASE__IS_RST_INVERTED    32'h0000000e
`define PLLE4_BASE__IS_RST_INVERTED_SZ 1

`define PLLE4_BASE__REF_JITTER    32'h0000000f
`define PLLE4_BASE__REF_JITTER_SZ 64

`define PLLE4_BASE__STARTUP_WAIT    32'h00000010
`define PLLE4_BASE__STARTUP_WAIT_SZ 40

`endif  // B_PLLE4_BASE_DEFINES_VH