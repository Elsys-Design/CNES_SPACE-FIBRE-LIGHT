// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_URAM288E5_DEFINES_VH
`else
`define B_URAM288E5_DEFINES_VH

// Look-up table parameters
//

`define URAM288E5_ADDR_N  1070
`define URAM288E5_ADDR_SZ 32
`define URAM288E5_DATA_SZ 288

// Attribute addresses
//

`define URAM288E5__AUTO_SLEEP_LATENCY    32'h00000000
`define URAM288E5__AUTO_SLEEP_LATENCY_SZ 32

`define URAM288E5__AVG_CONS_INACTIVE_CYCLES    32'h00000001
`define URAM288E5__AVG_CONS_INACTIVE_CYCLES_SZ 32

`define URAM288E5__BWE_MODE_A    32'h00000002
`define URAM288E5__BWE_MODE_A_SZ 144

`define URAM288E5__BWE_MODE_B    32'h00000003
`define URAM288E5__BWE_MODE_B_SZ 144

`define URAM288E5__CASCADE_ORDER_CTRL_A    32'h00000004
`define URAM288E5__CASCADE_ORDER_CTRL_A_SZ 48

`define URAM288E5__CASCADE_ORDER_CTRL_B    32'h00000005
`define URAM288E5__CASCADE_ORDER_CTRL_B_SZ 48

`define URAM288E5__CASCADE_ORDER_DATA_A    32'h00000006
`define URAM288E5__CASCADE_ORDER_DATA_A_SZ 48

`define URAM288E5__CASCADE_ORDER_DATA_B    32'h00000007
`define URAM288E5__CASCADE_ORDER_DATA_B_SZ 48

`define URAM288E5__EN_AUTO_SLEEP_MODE    32'h00000008
`define URAM288E5__EN_AUTO_SLEEP_MODE_SZ 40

`define URAM288E5__EN_ECC_RD_A    32'h00000009
`define URAM288E5__EN_ECC_RD_A_SZ 40

`define URAM288E5__EN_ECC_RD_B    32'h0000000a
`define URAM288E5__EN_ECC_RD_B_SZ 40

`define URAM288E5__EN_ECC_WR_A    32'h0000000b
`define URAM288E5__EN_ECC_WR_A_SZ 40

`define URAM288E5__EN_ECC_WR_B    32'h0000000c
`define URAM288E5__EN_ECC_WR_B_SZ 40

`define URAM288E5__INIT_000    32'h0000000d
`define URAM288E5__INIT_000_SZ 288

`define URAM288E5__INIT_001    32'h0000000e
`define URAM288E5__INIT_001_SZ 288

`define URAM288E5__INIT_002    32'h0000000f
`define URAM288E5__INIT_002_SZ 288

`define URAM288E5__INIT_003    32'h00000010
`define URAM288E5__INIT_003_SZ 288

`define URAM288E5__INIT_004    32'h00000011
`define URAM288E5__INIT_004_SZ 288

`define URAM288E5__INIT_005    32'h00000012
`define URAM288E5__INIT_005_SZ 288

`define URAM288E5__INIT_006    32'h00000013
`define URAM288E5__INIT_006_SZ 288

`define URAM288E5__INIT_007    32'h00000014
`define URAM288E5__INIT_007_SZ 288

`define URAM288E5__INIT_008    32'h00000015
`define URAM288E5__INIT_008_SZ 288

`define URAM288E5__INIT_009    32'h00000016
`define URAM288E5__INIT_009_SZ 288

`define URAM288E5__INIT_00A    32'h00000017
`define URAM288E5__INIT_00A_SZ 288

`define URAM288E5__INIT_00B    32'h00000018
`define URAM288E5__INIT_00B_SZ 288

`define URAM288E5__INIT_00C    32'h00000019
`define URAM288E5__INIT_00C_SZ 288

`define URAM288E5__INIT_00D    32'h0000001a
`define URAM288E5__INIT_00D_SZ 288

`define URAM288E5__INIT_00E    32'h0000001b
`define URAM288E5__INIT_00E_SZ 288

`define URAM288E5__INIT_00F    32'h0000001c
`define URAM288E5__INIT_00F_SZ 288

`define URAM288E5__INIT_010    32'h0000001d
`define URAM288E5__INIT_010_SZ 288

`define URAM288E5__INIT_011    32'h0000001e
`define URAM288E5__INIT_011_SZ 288

`define URAM288E5__INIT_012    32'h0000001f
`define URAM288E5__INIT_012_SZ 288

`define URAM288E5__INIT_013    32'h00000020
`define URAM288E5__INIT_013_SZ 288

`define URAM288E5__INIT_014    32'h00000021
`define URAM288E5__INIT_014_SZ 288

`define URAM288E5__INIT_015    32'h00000022
`define URAM288E5__INIT_015_SZ 288

`define URAM288E5__INIT_016    32'h00000023
`define URAM288E5__INIT_016_SZ 288

`define URAM288E5__INIT_017    32'h00000024
`define URAM288E5__INIT_017_SZ 288

`define URAM288E5__INIT_018    32'h00000025
`define URAM288E5__INIT_018_SZ 288

`define URAM288E5__INIT_019    32'h00000026
`define URAM288E5__INIT_019_SZ 288

`define URAM288E5__INIT_01A    32'h00000027
`define URAM288E5__INIT_01A_SZ 288

`define URAM288E5__INIT_01B    32'h00000028
`define URAM288E5__INIT_01B_SZ 288

`define URAM288E5__INIT_01C    32'h00000029
`define URAM288E5__INIT_01C_SZ 288

`define URAM288E5__INIT_01D    32'h0000002a
`define URAM288E5__INIT_01D_SZ 288

`define URAM288E5__INIT_01E    32'h0000002b
`define URAM288E5__INIT_01E_SZ 288

`define URAM288E5__INIT_01F    32'h0000002c
`define URAM288E5__INIT_01F_SZ 288

`define URAM288E5__INIT_020    32'h0000002d
`define URAM288E5__INIT_020_SZ 288

`define URAM288E5__INIT_021    32'h0000002e
`define URAM288E5__INIT_021_SZ 288

`define URAM288E5__INIT_022    32'h0000002f
`define URAM288E5__INIT_022_SZ 288

`define URAM288E5__INIT_023    32'h00000030
`define URAM288E5__INIT_023_SZ 288

`define URAM288E5__INIT_024    32'h00000031
`define URAM288E5__INIT_024_SZ 288

`define URAM288E5__INIT_025    32'h00000032
`define URAM288E5__INIT_025_SZ 288

`define URAM288E5__INIT_026    32'h00000033
`define URAM288E5__INIT_026_SZ 288

`define URAM288E5__INIT_027    32'h00000034
`define URAM288E5__INIT_027_SZ 288

`define URAM288E5__INIT_028    32'h00000035
`define URAM288E5__INIT_028_SZ 288

`define URAM288E5__INIT_029    32'h00000036
`define URAM288E5__INIT_029_SZ 288

`define URAM288E5__INIT_02A    32'h00000037
`define URAM288E5__INIT_02A_SZ 288

`define URAM288E5__INIT_02B    32'h00000038
`define URAM288E5__INIT_02B_SZ 288

`define URAM288E5__INIT_02C    32'h00000039
`define URAM288E5__INIT_02C_SZ 288

`define URAM288E5__INIT_02D    32'h0000003a
`define URAM288E5__INIT_02D_SZ 288

`define URAM288E5__INIT_02E    32'h0000003b
`define URAM288E5__INIT_02E_SZ 288

`define URAM288E5__INIT_02F    32'h0000003c
`define URAM288E5__INIT_02F_SZ 288

`define URAM288E5__INIT_030    32'h0000003d
`define URAM288E5__INIT_030_SZ 288

`define URAM288E5__INIT_031    32'h0000003e
`define URAM288E5__INIT_031_SZ 288

`define URAM288E5__INIT_032    32'h0000003f
`define URAM288E5__INIT_032_SZ 288

`define URAM288E5__INIT_033    32'h00000040
`define URAM288E5__INIT_033_SZ 288

`define URAM288E5__INIT_034    32'h00000041
`define URAM288E5__INIT_034_SZ 288

`define URAM288E5__INIT_035    32'h00000042
`define URAM288E5__INIT_035_SZ 288

`define URAM288E5__INIT_036    32'h00000043
`define URAM288E5__INIT_036_SZ 288

`define URAM288E5__INIT_037    32'h00000044
`define URAM288E5__INIT_037_SZ 288

`define URAM288E5__INIT_038    32'h00000045
`define URAM288E5__INIT_038_SZ 288

`define URAM288E5__INIT_039    32'h00000046
`define URAM288E5__INIT_039_SZ 288

`define URAM288E5__INIT_03A    32'h00000047
`define URAM288E5__INIT_03A_SZ 288

`define URAM288E5__INIT_03B    32'h00000048
`define URAM288E5__INIT_03B_SZ 288

`define URAM288E5__INIT_03C    32'h00000049
`define URAM288E5__INIT_03C_SZ 288

`define URAM288E5__INIT_03D    32'h0000004a
`define URAM288E5__INIT_03D_SZ 288

`define URAM288E5__INIT_03E    32'h0000004b
`define URAM288E5__INIT_03E_SZ 288

`define URAM288E5__INIT_03F    32'h0000004c
`define URAM288E5__INIT_03F_SZ 288

`define URAM288E5__INIT_040    32'h0000004d
`define URAM288E5__INIT_040_SZ 288

`define URAM288E5__INIT_041    32'h0000004e
`define URAM288E5__INIT_041_SZ 288

`define URAM288E5__INIT_042    32'h0000004f
`define URAM288E5__INIT_042_SZ 288

`define URAM288E5__INIT_043    32'h00000050
`define URAM288E5__INIT_043_SZ 288

`define URAM288E5__INIT_044    32'h00000051
`define URAM288E5__INIT_044_SZ 288

`define URAM288E5__INIT_045    32'h00000052
`define URAM288E5__INIT_045_SZ 288

`define URAM288E5__INIT_046    32'h00000053
`define URAM288E5__INIT_046_SZ 288

`define URAM288E5__INIT_047    32'h00000054
`define URAM288E5__INIT_047_SZ 288

`define URAM288E5__INIT_048    32'h00000055
`define URAM288E5__INIT_048_SZ 288

`define URAM288E5__INIT_049    32'h00000056
`define URAM288E5__INIT_049_SZ 288

`define URAM288E5__INIT_04A    32'h00000057
`define URAM288E5__INIT_04A_SZ 288

`define URAM288E5__INIT_04B    32'h00000058
`define URAM288E5__INIT_04B_SZ 288

`define URAM288E5__INIT_04C    32'h00000059
`define URAM288E5__INIT_04C_SZ 288

`define URAM288E5__INIT_04D    32'h0000005a
`define URAM288E5__INIT_04D_SZ 288

`define URAM288E5__INIT_04E    32'h0000005b
`define URAM288E5__INIT_04E_SZ 288

`define URAM288E5__INIT_04F    32'h0000005c
`define URAM288E5__INIT_04F_SZ 288

`define URAM288E5__INIT_050    32'h0000005d
`define URAM288E5__INIT_050_SZ 288

`define URAM288E5__INIT_051    32'h0000005e
`define URAM288E5__INIT_051_SZ 288

`define URAM288E5__INIT_052    32'h0000005f
`define URAM288E5__INIT_052_SZ 288

`define URAM288E5__INIT_053    32'h00000060
`define URAM288E5__INIT_053_SZ 288

`define URAM288E5__INIT_054    32'h00000061
`define URAM288E5__INIT_054_SZ 288

`define URAM288E5__INIT_055    32'h00000062
`define URAM288E5__INIT_055_SZ 288

`define URAM288E5__INIT_056    32'h00000063
`define URAM288E5__INIT_056_SZ 288

`define URAM288E5__INIT_057    32'h00000064
`define URAM288E5__INIT_057_SZ 288

`define URAM288E5__INIT_058    32'h00000065
`define URAM288E5__INIT_058_SZ 288

`define URAM288E5__INIT_059    32'h00000066
`define URAM288E5__INIT_059_SZ 288

`define URAM288E5__INIT_05A    32'h00000067
`define URAM288E5__INIT_05A_SZ 288

`define URAM288E5__INIT_05B    32'h00000068
`define URAM288E5__INIT_05B_SZ 288

`define URAM288E5__INIT_05C    32'h00000069
`define URAM288E5__INIT_05C_SZ 288

`define URAM288E5__INIT_05D    32'h0000006a
`define URAM288E5__INIT_05D_SZ 288

`define URAM288E5__INIT_05E    32'h0000006b
`define URAM288E5__INIT_05E_SZ 288

`define URAM288E5__INIT_05F    32'h0000006c
`define URAM288E5__INIT_05F_SZ 288

`define URAM288E5__INIT_060    32'h0000006d
`define URAM288E5__INIT_060_SZ 288

`define URAM288E5__INIT_061    32'h0000006e
`define URAM288E5__INIT_061_SZ 288

`define URAM288E5__INIT_062    32'h0000006f
`define URAM288E5__INIT_062_SZ 288

`define URAM288E5__INIT_063    32'h00000070
`define URAM288E5__INIT_063_SZ 288

`define URAM288E5__INIT_064    32'h00000071
`define URAM288E5__INIT_064_SZ 288

`define URAM288E5__INIT_065    32'h00000072
`define URAM288E5__INIT_065_SZ 288

`define URAM288E5__INIT_066    32'h00000073
`define URAM288E5__INIT_066_SZ 288

`define URAM288E5__INIT_067    32'h00000074
`define URAM288E5__INIT_067_SZ 288

`define URAM288E5__INIT_068    32'h00000075
`define URAM288E5__INIT_068_SZ 288

`define URAM288E5__INIT_069    32'h00000076
`define URAM288E5__INIT_069_SZ 288

`define URAM288E5__INIT_06A    32'h00000077
`define URAM288E5__INIT_06A_SZ 288

`define URAM288E5__INIT_06B    32'h00000078
`define URAM288E5__INIT_06B_SZ 288

`define URAM288E5__INIT_06C    32'h00000079
`define URAM288E5__INIT_06C_SZ 288

`define URAM288E5__INIT_06D    32'h0000007a
`define URAM288E5__INIT_06D_SZ 288

`define URAM288E5__INIT_06E    32'h0000007b
`define URAM288E5__INIT_06E_SZ 288

`define URAM288E5__INIT_06F    32'h0000007c
`define URAM288E5__INIT_06F_SZ 288

`define URAM288E5__INIT_070    32'h0000007d
`define URAM288E5__INIT_070_SZ 288

`define URAM288E5__INIT_071    32'h0000007e
`define URAM288E5__INIT_071_SZ 288

`define URAM288E5__INIT_072    32'h0000007f
`define URAM288E5__INIT_072_SZ 288

`define URAM288E5__INIT_073    32'h00000080
`define URAM288E5__INIT_073_SZ 288

`define URAM288E5__INIT_074    32'h00000081
`define URAM288E5__INIT_074_SZ 288

`define URAM288E5__INIT_075    32'h00000082
`define URAM288E5__INIT_075_SZ 288

`define URAM288E5__INIT_076    32'h00000083
`define URAM288E5__INIT_076_SZ 288

`define URAM288E5__INIT_077    32'h00000084
`define URAM288E5__INIT_077_SZ 288

`define URAM288E5__INIT_078    32'h00000085
`define URAM288E5__INIT_078_SZ 288

`define URAM288E5__INIT_079    32'h00000086
`define URAM288E5__INIT_079_SZ 288

`define URAM288E5__INIT_07A    32'h00000087
`define URAM288E5__INIT_07A_SZ 288

`define URAM288E5__INIT_07B    32'h00000088
`define URAM288E5__INIT_07B_SZ 288

`define URAM288E5__INIT_07C    32'h00000089
`define URAM288E5__INIT_07C_SZ 288

`define URAM288E5__INIT_07D    32'h0000008a
`define URAM288E5__INIT_07D_SZ 288

`define URAM288E5__INIT_07E    32'h0000008b
`define URAM288E5__INIT_07E_SZ 288

`define URAM288E5__INIT_07F    32'h0000008c
`define URAM288E5__INIT_07F_SZ 288

`define URAM288E5__INIT_080    32'h0000008d
`define URAM288E5__INIT_080_SZ 288

`define URAM288E5__INIT_081    32'h0000008e
`define URAM288E5__INIT_081_SZ 288

`define URAM288E5__INIT_082    32'h0000008f
`define URAM288E5__INIT_082_SZ 288

`define URAM288E5__INIT_083    32'h00000090
`define URAM288E5__INIT_083_SZ 288

`define URAM288E5__INIT_084    32'h00000091
`define URAM288E5__INIT_084_SZ 288

`define URAM288E5__INIT_085    32'h00000092
`define URAM288E5__INIT_085_SZ 288

`define URAM288E5__INIT_086    32'h00000093
`define URAM288E5__INIT_086_SZ 288

`define URAM288E5__INIT_087    32'h00000094
`define URAM288E5__INIT_087_SZ 288

`define URAM288E5__INIT_088    32'h00000095
`define URAM288E5__INIT_088_SZ 288

`define URAM288E5__INIT_089    32'h00000096
`define URAM288E5__INIT_089_SZ 288

`define URAM288E5__INIT_08A    32'h00000097
`define URAM288E5__INIT_08A_SZ 288

`define URAM288E5__INIT_08B    32'h00000098
`define URAM288E5__INIT_08B_SZ 288

`define URAM288E5__INIT_08C    32'h00000099
`define URAM288E5__INIT_08C_SZ 288

`define URAM288E5__INIT_08D    32'h0000009a
`define URAM288E5__INIT_08D_SZ 288

`define URAM288E5__INIT_08E    32'h0000009b
`define URAM288E5__INIT_08E_SZ 288

`define URAM288E5__INIT_08F    32'h0000009c
`define URAM288E5__INIT_08F_SZ 288

`define URAM288E5__INIT_090    32'h0000009d
`define URAM288E5__INIT_090_SZ 288

`define URAM288E5__INIT_091    32'h0000009e
`define URAM288E5__INIT_091_SZ 288

`define URAM288E5__INIT_092    32'h0000009f
`define URAM288E5__INIT_092_SZ 288

`define URAM288E5__INIT_093    32'h000000a0
`define URAM288E5__INIT_093_SZ 288

`define URAM288E5__INIT_094    32'h000000a1
`define URAM288E5__INIT_094_SZ 288

`define URAM288E5__INIT_095    32'h000000a2
`define URAM288E5__INIT_095_SZ 288

`define URAM288E5__INIT_096    32'h000000a3
`define URAM288E5__INIT_096_SZ 288

`define URAM288E5__INIT_097    32'h000000a4
`define URAM288E5__INIT_097_SZ 288

`define URAM288E5__INIT_098    32'h000000a5
`define URAM288E5__INIT_098_SZ 288

`define URAM288E5__INIT_099    32'h000000a6
`define URAM288E5__INIT_099_SZ 288

`define URAM288E5__INIT_09A    32'h000000a7
`define URAM288E5__INIT_09A_SZ 288

`define URAM288E5__INIT_09B    32'h000000a8
`define URAM288E5__INIT_09B_SZ 288

`define URAM288E5__INIT_09C    32'h000000a9
`define URAM288E5__INIT_09C_SZ 288

`define URAM288E5__INIT_09D    32'h000000aa
`define URAM288E5__INIT_09D_SZ 288

`define URAM288E5__INIT_09E    32'h000000ab
`define URAM288E5__INIT_09E_SZ 288

`define URAM288E5__INIT_09F    32'h000000ac
`define URAM288E5__INIT_09F_SZ 288

`define URAM288E5__INIT_0A0    32'h000000ad
`define URAM288E5__INIT_0A0_SZ 288

`define URAM288E5__INIT_0A1    32'h000000ae
`define URAM288E5__INIT_0A1_SZ 288

`define URAM288E5__INIT_0A2    32'h000000af
`define URAM288E5__INIT_0A2_SZ 288

`define URAM288E5__INIT_0A3    32'h000000b0
`define URAM288E5__INIT_0A3_SZ 288

`define URAM288E5__INIT_0A4    32'h000000b1
`define URAM288E5__INIT_0A4_SZ 288

`define URAM288E5__INIT_0A5    32'h000000b2
`define URAM288E5__INIT_0A5_SZ 288

`define URAM288E5__INIT_0A6    32'h000000b3
`define URAM288E5__INIT_0A6_SZ 288

`define URAM288E5__INIT_0A7    32'h000000b4
`define URAM288E5__INIT_0A7_SZ 288

`define URAM288E5__INIT_0A8    32'h000000b5
`define URAM288E5__INIT_0A8_SZ 288

`define URAM288E5__INIT_0A9    32'h000000b6
`define URAM288E5__INIT_0A9_SZ 288

`define URAM288E5__INIT_0AA    32'h000000b7
`define URAM288E5__INIT_0AA_SZ 288

`define URAM288E5__INIT_0AB    32'h000000b8
`define URAM288E5__INIT_0AB_SZ 288

`define URAM288E5__INIT_0AC    32'h000000b9
`define URAM288E5__INIT_0AC_SZ 288

`define URAM288E5__INIT_0AD    32'h000000ba
`define URAM288E5__INIT_0AD_SZ 288

`define URAM288E5__INIT_0AE    32'h000000bb
`define URAM288E5__INIT_0AE_SZ 288

`define URAM288E5__INIT_0AF    32'h000000bc
`define URAM288E5__INIT_0AF_SZ 288

`define URAM288E5__INIT_0B0    32'h000000bd
`define URAM288E5__INIT_0B0_SZ 288

`define URAM288E5__INIT_0B1    32'h000000be
`define URAM288E5__INIT_0B1_SZ 288

`define URAM288E5__INIT_0B2    32'h000000bf
`define URAM288E5__INIT_0B2_SZ 288

`define URAM288E5__INIT_0B3    32'h000000c0
`define URAM288E5__INIT_0B3_SZ 288

`define URAM288E5__INIT_0B4    32'h000000c1
`define URAM288E5__INIT_0B4_SZ 288

`define URAM288E5__INIT_0B5    32'h000000c2
`define URAM288E5__INIT_0B5_SZ 288

`define URAM288E5__INIT_0B6    32'h000000c3
`define URAM288E5__INIT_0B6_SZ 288

`define URAM288E5__INIT_0B7    32'h000000c4
`define URAM288E5__INIT_0B7_SZ 288

`define URAM288E5__INIT_0B8    32'h000000c5
`define URAM288E5__INIT_0B8_SZ 288

`define URAM288E5__INIT_0B9    32'h000000c6
`define URAM288E5__INIT_0B9_SZ 288

`define URAM288E5__INIT_0BA    32'h000000c7
`define URAM288E5__INIT_0BA_SZ 288

`define URAM288E5__INIT_0BB    32'h000000c8
`define URAM288E5__INIT_0BB_SZ 288

`define URAM288E5__INIT_0BC    32'h000000c9
`define URAM288E5__INIT_0BC_SZ 288

`define URAM288E5__INIT_0BD    32'h000000ca
`define URAM288E5__INIT_0BD_SZ 288

`define URAM288E5__INIT_0BE    32'h000000cb
`define URAM288E5__INIT_0BE_SZ 288

`define URAM288E5__INIT_0BF    32'h000000cc
`define URAM288E5__INIT_0BF_SZ 288

`define URAM288E5__INIT_0C0    32'h000000cd
`define URAM288E5__INIT_0C0_SZ 288

`define URAM288E5__INIT_0C1    32'h000000ce
`define URAM288E5__INIT_0C1_SZ 288

`define URAM288E5__INIT_0C2    32'h000000cf
`define URAM288E5__INIT_0C2_SZ 288

`define URAM288E5__INIT_0C3    32'h000000d0
`define URAM288E5__INIT_0C3_SZ 288

`define URAM288E5__INIT_0C4    32'h000000d1
`define URAM288E5__INIT_0C4_SZ 288

`define URAM288E5__INIT_0C5    32'h000000d2
`define URAM288E5__INIT_0C5_SZ 288

`define URAM288E5__INIT_0C6    32'h000000d3
`define URAM288E5__INIT_0C6_SZ 288

`define URAM288E5__INIT_0C7    32'h000000d4
`define URAM288E5__INIT_0C7_SZ 288

`define URAM288E5__INIT_0C8    32'h000000d5
`define URAM288E5__INIT_0C8_SZ 288

`define URAM288E5__INIT_0C9    32'h000000d6
`define URAM288E5__INIT_0C9_SZ 288

`define URAM288E5__INIT_0CA    32'h000000d7
`define URAM288E5__INIT_0CA_SZ 288

`define URAM288E5__INIT_0CB    32'h000000d8
`define URAM288E5__INIT_0CB_SZ 288

`define URAM288E5__INIT_0CC    32'h000000d9
`define URAM288E5__INIT_0CC_SZ 288

`define URAM288E5__INIT_0CD    32'h000000da
`define URAM288E5__INIT_0CD_SZ 288

`define URAM288E5__INIT_0CE    32'h000000db
`define URAM288E5__INIT_0CE_SZ 288

`define URAM288E5__INIT_0CF    32'h000000dc
`define URAM288E5__INIT_0CF_SZ 288

`define URAM288E5__INIT_0D0    32'h000000dd
`define URAM288E5__INIT_0D0_SZ 288

`define URAM288E5__INIT_0D1    32'h000000de
`define URAM288E5__INIT_0D1_SZ 288

`define URAM288E5__INIT_0D2    32'h000000df
`define URAM288E5__INIT_0D2_SZ 288

`define URAM288E5__INIT_0D3    32'h000000e0
`define URAM288E5__INIT_0D3_SZ 288

`define URAM288E5__INIT_0D4    32'h000000e1
`define URAM288E5__INIT_0D4_SZ 288

`define URAM288E5__INIT_0D5    32'h000000e2
`define URAM288E5__INIT_0D5_SZ 288

`define URAM288E5__INIT_0D6    32'h000000e3
`define URAM288E5__INIT_0D6_SZ 288

`define URAM288E5__INIT_0D7    32'h000000e4
`define URAM288E5__INIT_0D7_SZ 288

`define URAM288E5__INIT_0D8    32'h000000e5
`define URAM288E5__INIT_0D8_SZ 288

`define URAM288E5__INIT_0D9    32'h000000e6
`define URAM288E5__INIT_0D9_SZ 288

`define URAM288E5__INIT_0DA    32'h000000e7
`define URAM288E5__INIT_0DA_SZ 288

`define URAM288E5__INIT_0DB    32'h000000e8
`define URAM288E5__INIT_0DB_SZ 288

`define URAM288E5__INIT_0DC    32'h000000e9
`define URAM288E5__INIT_0DC_SZ 288

`define URAM288E5__INIT_0DD    32'h000000ea
`define URAM288E5__INIT_0DD_SZ 288

`define URAM288E5__INIT_0DE    32'h000000eb
`define URAM288E5__INIT_0DE_SZ 288

`define URAM288E5__INIT_0DF    32'h000000ec
`define URAM288E5__INIT_0DF_SZ 288

`define URAM288E5__INIT_0E0    32'h000000ed
`define URAM288E5__INIT_0E0_SZ 288

`define URAM288E5__INIT_0E1    32'h000000ee
`define URAM288E5__INIT_0E1_SZ 288

`define URAM288E5__INIT_0E2    32'h000000ef
`define URAM288E5__INIT_0E2_SZ 288

`define URAM288E5__INIT_0E3    32'h000000f0
`define URAM288E5__INIT_0E3_SZ 288

`define URAM288E5__INIT_0E4    32'h000000f1
`define URAM288E5__INIT_0E4_SZ 288

`define URAM288E5__INIT_0E5    32'h000000f2
`define URAM288E5__INIT_0E5_SZ 288

`define URAM288E5__INIT_0E6    32'h000000f3
`define URAM288E5__INIT_0E6_SZ 288

`define URAM288E5__INIT_0E7    32'h000000f4
`define URAM288E5__INIT_0E7_SZ 288

`define URAM288E5__INIT_0E8    32'h000000f5
`define URAM288E5__INIT_0E8_SZ 288

`define URAM288E5__INIT_0E9    32'h000000f6
`define URAM288E5__INIT_0E9_SZ 288

`define URAM288E5__INIT_0EA    32'h000000f7
`define URAM288E5__INIT_0EA_SZ 288

`define URAM288E5__INIT_0EB    32'h000000f8
`define URAM288E5__INIT_0EB_SZ 288

`define URAM288E5__INIT_0EC    32'h000000f9
`define URAM288E5__INIT_0EC_SZ 288

`define URAM288E5__INIT_0ED    32'h000000fa
`define URAM288E5__INIT_0ED_SZ 288

`define URAM288E5__INIT_0EE    32'h000000fb
`define URAM288E5__INIT_0EE_SZ 288

`define URAM288E5__INIT_0EF    32'h000000fc
`define URAM288E5__INIT_0EF_SZ 288

`define URAM288E5__INIT_0F0    32'h000000fd
`define URAM288E5__INIT_0F0_SZ 288

`define URAM288E5__INIT_0F1    32'h000000fe
`define URAM288E5__INIT_0F1_SZ 288

`define URAM288E5__INIT_0F2    32'h000000ff
`define URAM288E5__INIT_0F2_SZ 288

`define URAM288E5__INIT_0F3    32'h00000100
`define URAM288E5__INIT_0F3_SZ 288

`define URAM288E5__INIT_0F4    32'h00000101
`define URAM288E5__INIT_0F4_SZ 288

`define URAM288E5__INIT_0F5    32'h00000102
`define URAM288E5__INIT_0F5_SZ 288

`define URAM288E5__INIT_0F6    32'h00000103
`define URAM288E5__INIT_0F6_SZ 288

`define URAM288E5__INIT_0F7    32'h00000104
`define URAM288E5__INIT_0F7_SZ 288

`define URAM288E5__INIT_0F8    32'h00000105
`define URAM288E5__INIT_0F8_SZ 288

`define URAM288E5__INIT_0F9    32'h00000106
`define URAM288E5__INIT_0F9_SZ 288

`define URAM288E5__INIT_0FA    32'h00000107
`define URAM288E5__INIT_0FA_SZ 288

`define URAM288E5__INIT_0FB    32'h00000108
`define URAM288E5__INIT_0FB_SZ 288

`define URAM288E5__INIT_0FC    32'h00000109
`define URAM288E5__INIT_0FC_SZ 288

`define URAM288E5__INIT_0FD    32'h0000010a
`define URAM288E5__INIT_0FD_SZ 288

`define URAM288E5__INIT_0FE    32'h0000010b
`define URAM288E5__INIT_0FE_SZ 288

`define URAM288E5__INIT_0FF    32'h0000010c
`define URAM288E5__INIT_0FF_SZ 288

`define URAM288E5__INIT_100    32'h0000010d
`define URAM288E5__INIT_100_SZ 288

`define URAM288E5__INIT_101    32'h0000010e
`define URAM288E5__INIT_101_SZ 288

`define URAM288E5__INIT_102    32'h0000010f
`define URAM288E5__INIT_102_SZ 288

`define URAM288E5__INIT_103    32'h00000110
`define URAM288E5__INIT_103_SZ 288

`define URAM288E5__INIT_104    32'h00000111
`define URAM288E5__INIT_104_SZ 288

`define URAM288E5__INIT_105    32'h00000112
`define URAM288E5__INIT_105_SZ 288

`define URAM288E5__INIT_106    32'h00000113
`define URAM288E5__INIT_106_SZ 288

`define URAM288E5__INIT_107    32'h00000114
`define URAM288E5__INIT_107_SZ 288

`define URAM288E5__INIT_108    32'h00000115
`define URAM288E5__INIT_108_SZ 288

`define URAM288E5__INIT_109    32'h00000116
`define URAM288E5__INIT_109_SZ 288

`define URAM288E5__INIT_10A    32'h00000117
`define URAM288E5__INIT_10A_SZ 288

`define URAM288E5__INIT_10B    32'h00000118
`define URAM288E5__INIT_10B_SZ 288

`define URAM288E5__INIT_10C    32'h00000119
`define URAM288E5__INIT_10C_SZ 288

`define URAM288E5__INIT_10D    32'h0000011a
`define URAM288E5__INIT_10D_SZ 288

`define URAM288E5__INIT_10E    32'h0000011b
`define URAM288E5__INIT_10E_SZ 288

`define URAM288E5__INIT_10F    32'h0000011c
`define URAM288E5__INIT_10F_SZ 288

`define URAM288E5__INIT_110    32'h0000011d
`define URAM288E5__INIT_110_SZ 288

`define URAM288E5__INIT_111    32'h0000011e
`define URAM288E5__INIT_111_SZ 288

`define URAM288E5__INIT_112    32'h0000011f
`define URAM288E5__INIT_112_SZ 288

`define URAM288E5__INIT_113    32'h00000120
`define URAM288E5__INIT_113_SZ 288

`define URAM288E5__INIT_114    32'h00000121
`define URAM288E5__INIT_114_SZ 288

`define URAM288E5__INIT_115    32'h00000122
`define URAM288E5__INIT_115_SZ 288

`define URAM288E5__INIT_116    32'h00000123
`define URAM288E5__INIT_116_SZ 288

`define URAM288E5__INIT_117    32'h00000124
`define URAM288E5__INIT_117_SZ 288

`define URAM288E5__INIT_118    32'h00000125
`define URAM288E5__INIT_118_SZ 288

`define URAM288E5__INIT_119    32'h00000126
`define URAM288E5__INIT_119_SZ 288

`define URAM288E5__INIT_11A    32'h00000127
`define URAM288E5__INIT_11A_SZ 288

`define URAM288E5__INIT_11B    32'h00000128
`define URAM288E5__INIT_11B_SZ 288

`define URAM288E5__INIT_11C    32'h00000129
`define URAM288E5__INIT_11C_SZ 288

`define URAM288E5__INIT_11D    32'h0000012a
`define URAM288E5__INIT_11D_SZ 288

`define URAM288E5__INIT_11E    32'h0000012b
`define URAM288E5__INIT_11E_SZ 288

`define URAM288E5__INIT_11F    32'h0000012c
`define URAM288E5__INIT_11F_SZ 288

`define URAM288E5__INIT_120    32'h0000012d
`define URAM288E5__INIT_120_SZ 288

`define URAM288E5__INIT_121    32'h0000012e
`define URAM288E5__INIT_121_SZ 288

`define URAM288E5__INIT_122    32'h0000012f
`define URAM288E5__INIT_122_SZ 288

`define URAM288E5__INIT_123    32'h00000130
`define URAM288E5__INIT_123_SZ 288

`define URAM288E5__INIT_124    32'h00000131
`define URAM288E5__INIT_124_SZ 288

`define URAM288E5__INIT_125    32'h00000132
`define URAM288E5__INIT_125_SZ 288

`define URAM288E5__INIT_126    32'h00000133
`define URAM288E5__INIT_126_SZ 288

`define URAM288E5__INIT_127    32'h00000134
`define URAM288E5__INIT_127_SZ 288

`define URAM288E5__INIT_128    32'h00000135
`define URAM288E5__INIT_128_SZ 288

`define URAM288E5__INIT_129    32'h00000136
`define URAM288E5__INIT_129_SZ 288

`define URAM288E5__INIT_12A    32'h00000137
`define URAM288E5__INIT_12A_SZ 288

`define URAM288E5__INIT_12B    32'h00000138
`define URAM288E5__INIT_12B_SZ 288

`define URAM288E5__INIT_12C    32'h00000139
`define URAM288E5__INIT_12C_SZ 288

`define URAM288E5__INIT_12D    32'h0000013a
`define URAM288E5__INIT_12D_SZ 288

`define URAM288E5__INIT_12E    32'h0000013b
`define URAM288E5__INIT_12E_SZ 288

`define URAM288E5__INIT_12F    32'h0000013c
`define URAM288E5__INIT_12F_SZ 288

`define URAM288E5__INIT_130    32'h0000013d
`define URAM288E5__INIT_130_SZ 288

`define URAM288E5__INIT_131    32'h0000013e
`define URAM288E5__INIT_131_SZ 288

`define URAM288E5__INIT_132    32'h0000013f
`define URAM288E5__INIT_132_SZ 288

`define URAM288E5__INIT_133    32'h00000140
`define URAM288E5__INIT_133_SZ 288

`define URAM288E5__INIT_134    32'h00000141
`define URAM288E5__INIT_134_SZ 288

`define URAM288E5__INIT_135    32'h00000142
`define URAM288E5__INIT_135_SZ 288

`define URAM288E5__INIT_136    32'h00000143
`define URAM288E5__INIT_136_SZ 288

`define URAM288E5__INIT_137    32'h00000144
`define URAM288E5__INIT_137_SZ 288

`define URAM288E5__INIT_138    32'h00000145
`define URAM288E5__INIT_138_SZ 288

`define URAM288E5__INIT_139    32'h00000146
`define URAM288E5__INIT_139_SZ 288

`define URAM288E5__INIT_13A    32'h00000147
`define URAM288E5__INIT_13A_SZ 288

`define URAM288E5__INIT_13B    32'h00000148
`define URAM288E5__INIT_13B_SZ 288

`define URAM288E5__INIT_13C    32'h00000149
`define URAM288E5__INIT_13C_SZ 288

`define URAM288E5__INIT_13D    32'h0000014a
`define URAM288E5__INIT_13D_SZ 288

`define URAM288E5__INIT_13E    32'h0000014b
`define URAM288E5__INIT_13E_SZ 288

`define URAM288E5__INIT_13F    32'h0000014c
`define URAM288E5__INIT_13F_SZ 288

`define URAM288E5__INIT_140    32'h0000014d
`define URAM288E5__INIT_140_SZ 288

`define URAM288E5__INIT_141    32'h0000014e
`define URAM288E5__INIT_141_SZ 288

`define URAM288E5__INIT_142    32'h0000014f
`define URAM288E5__INIT_142_SZ 288

`define URAM288E5__INIT_143    32'h00000150
`define URAM288E5__INIT_143_SZ 288

`define URAM288E5__INIT_144    32'h00000151
`define URAM288E5__INIT_144_SZ 288

`define URAM288E5__INIT_145    32'h00000152
`define URAM288E5__INIT_145_SZ 288

`define URAM288E5__INIT_146    32'h00000153
`define URAM288E5__INIT_146_SZ 288

`define URAM288E5__INIT_147    32'h00000154
`define URAM288E5__INIT_147_SZ 288

`define URAM288E5__INIT_148    32'h00000155
`define URAM288E5__INIT_148_SZ 288

`define URAM288E5__INIT_149    32'h00000156
`define URAM288E5__INIT_149_SZ 288

`define URAM288E5__INIT_14A    32'h00000157
`define URAM288E5__INIT_14A_SZ 288

`define URAM288E5__INIT_14B    32'h00000158
`define URAM288E5__INIT_14B_SZ 288

`define URAM288E5__INIT_14C    32'h00000159
`define URAM288E5__INIT_14C_SZ 288

`define URAM288E5__INIT_14D    32'h0000015a
`define URAM288E5__INIT_14D_SZ 288

`define URAM288E5__INIT_14E    32'h0000015b
`define URAM288E5__INIT_14E_SZ 288

`define URAM288E5__INIT_14F    32'h0000015c
`define URAM288E5__INIT_14F_SZ 288

`define URAM288E5__INIT_150    32'h0000015d
`define URAM288E5__INIT_150_SZ 288

`define URAM288E5__INIT_151    32'h0000015e
`define URAM288E5__INIT_151_SZ 288

`define URAM288E5__INIT_152    32'h0000015f
`define URAM288E5__INIT_152_SZ 288

`define URAM288E5__INIT_153    32'h00000160
`define URAM288E5__INIT_153_SZ 288

`define URAM288E5__INIT_154    32'h00000161
`define URAM288E5__INIT_154_SZ 288

`define URAM288E5__INIT_155    32'h00000162
`define URAM288E5__INIT_155_SZ 288

`define URAM288E5__INIT_156    32'h00000163
`define URAM288E5__INIT_156_SZ 288

`define URAM288E5__INIT_157    32'h00000164
`define URAM288E5__INIT_157_SZ 288

`define URAM288E5__INIT_158    32'h00000165
`define URAM288E5__INIT_158_SZ 288

`define URAM288E5__INIT_159    32'h00000166
`define URAM288E5__INIT_159_SZ 288

`define URAM288E5__INIT_15A    32'h00000167
`define URAM288E5__INIT_15A_SZ 288

`define URAM288E5__INIT_15B    32'h00000168
`define URAM288E5__INIT_15B_SZ 288

`define URAM288E5__INIT_15C    32'h00000169
`define URAM288E5__INIT_15C_SZ 288

`define URAM288E5__INIT_15D    32'h0000016a
`define URAM288E5__INIT_15D_SZ 288

`define URAM288E5__INIT_15E    32'h0000016b
`define URAM288E5__INIT_15E_SZ 288

`define URAM288E5__INIT_15F    32'h0000016c
`define URAM288E5__INIT_15F_SZ 288

`define URAM288E5__INIT_160    32'h0000016d
`define URAM288E5__INIT_160_SZ 288

`define URAM288E5__INIT_161    32'h0000016e
`define URAM288E5__INIT_161_SZ 288

`define URAM288E5__INIT_162    32'h0000016f
`define URAM288E5__INIT_162_SZ 288

`define URAM288E5__INIT_163    32'h00000170
`define URAM288E5__INIT_163_SZ 288

`define URAM288E5__INIT_164    32'h00000171
`define URAM288E5__INIT_164_SZ 288

`define URAM288E5__INIT_165    32'h00000172
`define URAM288E5__INIT_165_SZ 288

`define URAM288E5__INIT_166    32'h00000173
`define URAM288E5__INIT_166_SZ 288

`define URAM288E5__INIT_167    32'h00000174
`define URAM288E5__INIT_167_SZ 288

`define URAM288E5__INIT_168    32'h00000175
`define URAM288E5__INIT_168_SZ 288

`define URAM288E5__INIT_169    32'h00000176
`define URAM288E5__INIT_169_SZ 288

`define URAM288E5__INIT_16A    32'h00000177
`define URAM288E5__INIT_16A_SZ 288

`define URAM288E5__INIT_16B    32'h00000178
`define URAM288E5__INIT_16B_SZ 288

`define URAM288E5__INIT_16C    32'h00000179
`define URAM288E5__INIT_16C_SZ 288

`define URAM288E5__INIT_16D    32'h0000017a
`define URAM288E5__INIT_16D_SZ 288

`define URAM288E5__INIT_16E    32'h0000017b
`define URAM288E5__INIT_16E_SZ 288

`define URAM288E5__INIT_16F    32'h0000017c
`define URAM288E5__INIT_16F_SZ 288

`define URAM288E5__INIT_170    32'h0000017d
`define URAM288E5__INIT_170_SZ 288

`define URAM288E5__INIT_171    32'h0000017e
`define URAM288E5__INIT_171_SZ 288

`define URAM288E5__INIT_172    32'h0000017f
`define URAM288E5__INIT_172_SZ 288

`define URAM288E5__INIT_173    32'h00000180
`define URAM288E5__INIT_173_SZ 288

`define URAM288E5__INIT_174    32'h00000181
`define URAM288E5__INIT_174_SZ 288

`define URAM288E5__INIT_175    32'h00000182
`define URAM288E5__INIT_175_SZ 288

`define URAM288E5__INIT_176    32'h00000183
`define URAM288E5__INIT_176_SZ 288

`define URAM288E5__INIT_177    32'h00000184
`define URAM288E5__INIT_177_SZ 288

`define URAM288E5__INIT_178    32'h00000185
`define URAM288E5__INIT_178_SZ 288

`define URAM288E5__INIT_179    32'h00000186
`define URAM288E5__INIT_179_SZ 288

`define URAM288E5__INIT_17A    32'h00000187
`define URAM288E5__INIT_17A_SZ 288

`define URAM288E5__INIT_17B    32'h00000188
`define URAM288E5__INIT_17B_SZ 288

`define URAM288E5__INIT_17C    32'h00000189
`define URAM288E5__INIT_17C_SZ 288

`define URAM288E5__INIT_17D    32'h0000018a
`define URAM288E5__INIT_17D_SZ 288

`define URAM288E5__INIT_17E    32'h0000018b
`define URAM288E5__INIT_17E_SZ 288

`define URAM288E5__INIT_17F    32'h0000018c
`define URAM288E5__INIT_17F_SZ 288

`define URAM288E5__INIT_180    32'h0000018d
`define URAM288E5__INIT_180_SZ 288

`define URAM288E5__INIT_181    32'h0000018e
`define URAM288E5__INIT_181_SZ 288

`define URAM288E5__INIT_182    32'h0000018f
`define URAM288E5__INIT_182_SZ 288

`define URAM288E5__INIT_183    32'h00000190
`define URAM288E5__INIT_183_SZ 288

`define URAM288E5__INIT_184    32'h00000191
`define URAM288E5__INIT_184_SZ 288

`define URAM288E5__INIT_185    32'h00000192
`define URAM288E5__INIT_185_SZ 288

`define URAM288E5__INIT_186    32'h00000193
`define URAM288E5__INIT_186_SZ 288

`define URAM288E5__INIT_187    32'h00000194
`define URAM288E5__INIT_187_SZ 288

`define URAM288E5__INIT_188    32'h00000195
`define URAM288E5__INIT_188_SZ 288

`define URAM288E5__INIT_189    32'h00000196
`define URAM288E5__INIT_189_SZ 288

`define URAM288E5__INIT_18A    32'h00000197
`define URAM288E5__INIT_18A_SZ 288

`define URAM288E5__INIT_18B    32'h00000198
`define URAM288E5__INIT_18B_SZ 288

`define URAM288E5__INIT_18C    32'h00000199
`define URAM288E5__INIT_18C_SZ 288

`define URAM288E5__INIT_18D    32'h0000019a
`define URAM288E5__INIT_18D_SZ 288

`define URAM288E5__INIT_18E    32'h0000019b
`define URAM288E5__INIT_18E_SZ 288

`define URAM288E5__INIT_18F    32'h0000019c
`define URAM288E5__INIT_18F_SZ 288

`define URAM288E5__INIT_190    32'h0000019d
`define URAM288E5__INIT_190_SZ 288

`define URAM288E5__INIT_191    32'h0000019e
`define URAM288E5__INIT_191_SZ 288

`define URAM288E5__INIT_192    32'h0000019f
`define URAM288E5__INIT_192_SZ 288

`define URAM288E5__INIT_193    32'h000001a0
`define URAM288E5__INIT_193_SZ 288

`define URAM288E5__INIT_194    32'h000001a1
`define URAM288E5__INIT_194_SZ 288

`define URAM288E5__INIT_195    32'h000001a2
`define URAM288E5__INIT_195_SZ 288

`define URAM288E5__INIT_196    32'h000001a3
`define URAM288E5__INIT_196_SZ 288

`define URAM288E5__INIT_197    32'h000001a4
`define URAM288E5__INIT_197_SZ 288

`define URAM288E5__INIT_198    32'h000001a5
`define URAM288E5__INIT_198_SZ 288

`define URAM288E5__INIT_199    32'h000001a6
`define URAM288E5__INIT_199_SZ 288

`define URAM288E5__INIT_19A    32'h000001a7
`define URAM288E5__INIT_19A_SZ 288

`define URAM288E5__INIT_19B    32'h000001a8
`define URAM288E5__INIT_19B_SZ 288

`define URAM288E5__INIT_19C    32'h000001a9
`define URAM288E5__INIT_19C_SZ 288

`define URAM288E5__INIT_19D    32'h000001aa
`define URAM288E5__INIT_19D_SZ 288

`define URAM288E5__INIT_19E    32'h000001ab
`define URAM288E5__INIT_19E_SZ 288

`define URAM288E5__INIT_19F    32'h000001ac
`define URAM288E5__INIT_19F_SZ 288

`define URAM288E5__INIT_1A0    32'h000001ad
`define URAM288E5__INIT_1A0_SZ 288

`define URAM288E5__INIT_1A1    32'h000001ae
`define URAM288E5__INIT_1A1_SZ 288

`define URAM288E5__INIT_1A2    32'h000001af
`define URAM288E5__INIT_1A2_SZ 288

`define URAM288E5__INIT_1A3    32'h000001b0
`define URAM288E5__INIT_1A3_SZ 288

`define URAM288E5__INIT_1A4    32'h000001b1
`define URAM288E5__INIT_1A4_SZ 288

`define URAM288E5__INIT_1A5    32'h000001b2
`define URAM288E5__INIT_1A5_SZ 288

`define URAM288E5__INIT_1A6    32'h000001b3
`define URAM288E5__INIT_1A6_SZ 288

`define URAM288E5__INIT_1A7    32'h000001b4
`define URAM288E5__INIT_1A7_SZ 288

`define URAM288E5__INIT_1A8    32'h000001b5
`define URAM288E5__INIT_1A8_SZ 288

`define URAM288E5__INIT_1A9    32'h000001b6
`define URAM288E5__INIT_1A9_SZ 288

`define URAM288E5__INIT_1AA    32'h000001b7
`define URAM288E5__INIT_1AA_SZ 288

`define URAM288E5__INIT_1AB    32'h000001b8
`define URAM288E5__INIT_1AB_SZ 288

`define URAM288E5__INIT_1AC    32'h000001b9
`define URAM288E5__INIT_1AC_SZ 288

`define URAM288E5__INIT_1AD    32'h000001ba
`define URAM288E5__INIT_1AD_SZ 288

`define URAM288E5__INIT_1AE    32'h000001bb
`define URAM288E5__INIT_1AE_SZ 288

`define URAM288E5__INIT_1AF    32'h000001bc
`define URAM288E5__INIT_1AF_SZ 288

`define URAM288E5__INIT_1B0    32'h000001bd
`define URAM288E5__INIT_1B0_SZ 288

`define URAM288E5__INIT_1B1    32'h000001be
`define URAM288E5__INIT_1B1_SZ 288

`define URAM288E5__INIT_1B2    32'h000001bf
`define URAM288E5__INIT_1B2_SZ 288

`define URAM288E5__INIT_1B3    32'h000001c0
`define URAM288E5__INIT_1B3_SZ 288

`define URAM288E5__INIT_1B4    32'h000001c1
`define URAM288E5__INIT_1B4_SZ 288

`define URAM288E5__INIT_1B5    32'h000001c2
`define URAM288E5__INIT_1B5_SZ 288

`define URAM288E5__INIT_1B6    32'h000001c3
`define URAM288E5__INIT_1B6_SZ 288

`define URAM288E5__INIT_1B7    32'h000001c4
`define URAM288E5__INIT_1B7_SZ 288

`define URAM288E5__INIT_1B8    32'h000001c5
`define URAM288E5__INIT_1B8_SZ 288

`define URAM288E5__INIT_1B9    32'h000001c6
`define URAM288E5__INIT_1B9_SZ 288

`define URAM288E5__INIT_1BA    32'h000001c7
`define URAM288E5__INIT_1BA_SZ 288

`define URAM288E5__INIT_1BB    32'h000001c8
`define URAM288E5__INIT_1BB_SZ 288

`define URAM288E5__INIT_1BC    32'h000001c9
`define URAM288E5__INIT_1BC_SZ 288

`define URAM288E5__INIT_1BD    32'h000001ca
`define URAM288E5__INIT_1BD_SZ 288

`define URAM288E5__INIT_1BE    32'h000001cb
`define URAM288E5__INIT_1BE_SZ 288

`define URAM288E5__INIT_1BF    32'h000001cc
`define URAM288E5__INIT_1BF_SZ 288

`define URAM288E5__INIT_1C0    32'h000001cd
`define URAM288E5__INIT_1C0_SZ 288

`define URAM288E5__INIT_1C1    32'h000001ce
`define URAM288E5__INIT_1C1_SZ 288

`define URAM288E5__INIT_1C2    32'h000001cf
`define URAM288E5__INIT_1C2_SZ 288

`define URAM288E5__INIT_1C3    32'h000001d0
`define URAM288E5__INIT_1C3_SZ 288

`define URAM288E5__INIT_1C4    32'h000001d1
`define URAM288E5__INIT_1C4_SZ 288

`define URAM288E5__INIT_1C5    32'h000001d2
`define URAM288E5__INIT_1C5_SZ 288

`define URAM288E5__INIT_1C6    32'h000001d3
`define URAM288E5__INIT_1C6_SZ 288

`define URAM288E5__INIT_1C7    32'h000001d4
`define URAM288E5__INIT_1C7_SZ 288

`define URAM288E5__INIT_1C8    32'h000001d5
`define URAM288E5__INIT_1C8_SZ 288

`define URAM288E5__INIT_1C9    32'h000001d6
`define URAM288E5__INIT_1C9_SZ 288

`define URAM288E5__INIT_1CA    32'h000001d7
`define URAM288E5__INIT_1CA_SZ 288

`define URAM288E5__INIT_1CB    32'h000001d8
`define URAM288E5__INIT_1CB_SZ 288

`define URAM288E5__INIT_1CC    32'h000001d9
`define URAM288E5__INIT_1CC_SZ 288

`define URAM288E5__INIT_1CD    32'h000001da
`define URAM288E5__INIT_1CD_SZ 288

`define URAM288E5__INIT_1CE    32'h000001db
`define URAM288E5__INIT_1CE_SZ 288

`define URAM288E5__INIT_1CF    32'h000001dc
`define URAM288E5__INIT_1CF_SZ 288

`define URAM288E5__INIT_1D0    32'h000001dd
`define URAM288E5__INIT_1D0_SZ 288

`define URAM288E5__INIT_1D1    32'h000001de
`define URAM288E5__INIT_1D1_SZ 288

`define URAM288E5__INIT_1D2    32'h000001df
`define URAM288E5__INIT_1D2_SZ 288

`define URAM288E5__INIT_1D3    32'h000001e0
`define URAM288E5__INIT_1D3_SZ 288

`define URAM288E5__INIT_1D4    32'h000001e1
`define URAM288E5__INIT_1D4_SZ 288

`define URAM288E5__INIT_1D5    32'h000001e2
`define URAM288E5__INIT_1D5_SZ 288

`define URAM288E5__INIT_1D6    32'h000001e3
`define URAM288E5__INIT_1D6_SZ 288

`define URAM288E5__INIT_1D7    32'h000001e4
`define URAM288E5__INIT_1D7_SZ 288

`define URAM288E5__INIT_1D8    32'h000001e5
`define URAM288E5__INIT_1D8_SZ 288

`define URAM288E5__INIT_1D9    32'h000001e6
`define URAM288E5__INIT_1D9_SZ 288

`define URAM288E5__INIT_1DA    32'h000001e7
`define URAM288E5__INIT_1DA_SZ 288

`define URAM288E5__INIT_1DB    32'h000001e8
`define URAM288E5__INIT_1DB_SZ 288

`define URAM288E5__INIT_1DC    32'h000001e9
`define URAM288E5__INIT_1DC_SZ 288

`define URAM288E5__INIT_1DD    32'h000001ea
`define URAM288E5__INIT_1DD_SZ 288

`define URAM288E5__INIT_1DE    32'h000001eb
`define URAM288E5__INIT_1DE_SZ 288

`define URAM288E5__INIT_1DF    32'h000001ec
`define URAM288E5__INIT_1DF_SZ 288

`define URAM288E5__INIT_1E0    32'h000001ed
`define URAM288E5__INIT_1E0_SZ 288

`define URAM288E5__INIT_1E1    32'h000001ee
`define URAM288E5__INIT_1E1_SZ 288

`define URAM288E5__INIT_1E2    32'h000001ef
`define URAM288E5__INIT_1E2_SZ 288

`define URAM288E5__INIT_1E3    32'h000001f0
`define URAM288E5__INIT_1E3_SZ 288

`define URAM288E5__INIT_1E4    32'h000001f1
`define URAM288E5__INIT_1E4_SZ 288

`define URAM288E5__INIT_1E5    32'h000001f2
`define URAM288E5__INIT_1E5_SZ 288

`define URAM288E5__INIT_1E6    32'h000001f3
`define URAM288E5__INIT_1E6_SZ 288

`define URAM288E5__INIT_1E7    32'h000001f4
`define URAM288E5__INIT_1E7_SZ 288

`define URAM288E5__INIT_1E8    32'h000001f5
`define URAM288E5__INIT_1E8_SZ 288

`define URAM288E5__INIT_1E9    32'h000001f6
`define URAM288E5__INIT_1E9_SZ 288

`define URAM288E5__INIT_1EA    32'h000001f7
`define URAM288E5__INIT_1EA_SZ 288

`define URAM288E5__INIT_1EB    32'h000001f8
`define URAM288E5__INIT_1EB_SZ 288

`define URAM288E5__INIT_1EC    32'h000001f9
`define URAM288E5__INIT_1EC_SZ 288

`define URAM288E5__INIT_1ED    32'h000001fa
`define URAM288E5__INIT_1ED_SZ 288

`define URAM288E5__INIT_1EE    32'h000001fb
`define URAM288E5__INIT_1EE_SZ 288

`define URAM288E5__INIT_1EF    32'h000001fc
`define URAM288E5__INIT_1EF_SZ 288

`define URAM288E5__INIT_1F0    32'h000001fd
`define URAM288E5__INIT_1F0_SZ 288

`define URAM288E5__INIT_1F1    32'h000001fe
`define URAM288E5__INIT_1F1_SZ 288

`define URAM288E5__INIT_1F2    32'h000001ff
`define URAM288E5__INIT_1F2_SZ 288

`define URAM288E5__INIT_1F3    32'h00000200
`define URAM288E5__INIT_1F3_SZ 288

`define URAM288E5__INIT_1F4    32'h00000201
`define URAM288E5__INIT_1F4_SZ 288

`define URAM288E5__INIT_1F5    32'h00000202
`define URAM288E5__INIT_1F5_SZ 288

`define URAM288E5__INIT_1F6    32'h00000203
`define URAM288E5__INIT_1F6_SZ 288

`define URAM288E5__INIT_1F7    32'h00000204
`define URAM288E5__INIT_1F7_SZ 288

`define URAM288E5__INIT_1F8    32'h00000205
`define URAM288E5__INIT_1F8_SZ 288

`define URAM288E5__INIT_1F9    32'h00000206
`define URAM288E5__INIT_1F9_SZ 288

`define URAM288E5__INIT_1FA    32'h00000207
`define URAM288E5__INIT_1FA_SZ 288

`define URAM288E5__INIT_1FB    32'h00000208
`define URAM288E5__INIT_1FB_SZ 288

`define URAM288E5__INIT_1FC    32'h00000209
`define URAM288E5__INIT_1FC_SZ 288

`define URAM288E5__INIT_1FD    32'h0000020a
`define URAM288E5__INIT_1FD_SZ 288

`define URAM288E5__INIT_1FE    32'h0000020b
`define URAM288E5__INIT_1FE_SZ 288

`define URAM288E5__INIT_1FF    32'h0000020c
`define URAM288E5__INIT_1FF_SZ 288

`define URAM288E5__INIT_200    32'h0000020d
`define URAM288E5__INIT_200_SZ 288

`define URAM288E5__INIT_201    32'h0000020e
`define URAM288E5__INIT_201_SZ 288

`define URAM288E5__INIT_202    32'h0000020f
`define URAM288E5__INIT_202_SZ 288

`define URAM288E5__INIT_203    32'h00000210
`define URAM288E5__INIT_203_SZ 288

`define URAM288E5__INIT_204    32'h00000211
`define URAM288E5__INIT_204_SZ 288

`define URAM288E5__INIT_205    32'h00000212
`define URAM288E5__INIT_205_SZ 288

`define URAM288E5__INIT_206    32'h00000213
`define URAM288E5__INIT_206_SZ 288

`define URAM288E5__INIT_207    32'h00000214
`define URAM288E5__INIT_207_SZ 288

`define URAM288E5__INIT_208    32'h00000215
`define URAM288E5__INIT_208_SZ 288

`define URAM288E5__INIT_209    32'h00000216
`define URAM288E5__INIT_209_SZ 288

`define URAM288E5__INIT_20A    32'h00000217
`define URAM288E5__INIT_20A_SZ 288

`define URAM288E5__INIT_20B    32'h00000218
`define URAM288E5__INIT_20B_SZ 288

`define URAM288E5__INIT_20C    32'h00000219
`define URAM288E5__INIT_20C_SZ 288

`define URAM288E5__INIT_20D    32'h0000021a
`define URAM288E5__INIT_20D_SZ 288

`define URAM288E5__INIT_20E    32'h0000021b
`define URAM288E5__INIT_20E_SZ 288

`define URAM288E5__INIT_20F    32'h0000021c
`define URAM288E5__INIT_20F_SZ 288

`define URAM288E5__INIT_210    32'h0000021d
`define URAM288E5__INIT_210_SZ 288

`define URAM288E5__INIT_211    32'h0000021e
`define URAM288E5__INIT_211_SZ 288

`define URAM288E5__INIT_212    32'h0000021f
`define URAM288E5__INIT_212_SZ 288

`define URAM288E5__INIT_213    32'h00000220
`define URAM288E5__INIT_213_SZ 288

`define URAM288E5__INIT_214    32'h00000221
`define URAM288E5__INIT_214_SZ 288

`define URAM288E5__INIT_215    32'h00000222
`define URAM288E5__INIT_215_SZ 288

`define URAM288E5__INIT_216    32'h00000223
`define URAM288E5__INIT_216_SZ 288

`define URAM288E5__INIT_217    32'h00000224
`define URAM288E5__INIT_217_SZ 288

`define URAM288E5__INIT_218    32'h00000225
`define URAM288E5__INIT_218_SZ 288

`define URAM288E5__INIT_219    32'h00000226
`define URAM288E5__INIT_219_SZ 288

`define URAM288E5__INIT_21A    32'h00000227
`define URAM288E5__INIT_21A_SZ 288

`define URAM288E5__INIT_21B    32'h00000228
`define URAM288E5__INIT_21B_SZ 288

`define URAM288E5__INIT_21C    32'h00000229
`define URAM288E5__INIT_21C_SZ 288

`define URAM288E5__INIT_21D    32'h0000022a
`define URAM288E5__INIT_21D_SZ 288

`define URAM288E5__INIT_21E    32'h0000022b
`define URAM288E5__INIT_21E_SZ 288

`define URAM288E5__INIT_21F    32'h0000022c
`define URAM288E5__INIT_21F_SZ 288

`define URAM288E5__INIT_220    32'h0000022d
`define URAM288E5__INIT_220_SZ 288

`define URAM288E5__INIT_221    32'h0000022e
`define URAM288E5__INIT_221_SZ 288

`define URAM288E5__INIT_222    32'h0000022f
`define URAM288E5__INIT_222_SZ 288

`define URAM288E5__INIT_223    32'h00000230
`define URAM288E5__INIT_223_SZ 288

`define URAM288E5__INIT_224    32'h00000231
`define URAM288E5__INIT_224_SZ 288

`define URAM288E5__INIT_225    32'h00000232
`define URAM288E5__INIT_225_SZ 288

`define URAM288E5__INIT_226    32'h00000233
`define URAM288E5__INIT_226_SZ 288

`define URAM288E5__INIT_227    32'h00000234
`define URAM288E5__INIT_227_SZ 288

`define URAM288E5__INIT_228    32'h00000235
`define URAM288E5__INIT_228_SZ 288

`define URAM288E5__INIT_229    32'h00000236
`define URAM288E5__INIT_229_SZ 288

`define URAM288E5__INIT_22A    32'h00000237
`define URAM288E5__INIT_22A_SZ 288

`define URAM288E5__INIT_22B    32'h00000238
`define URAM288E5__INIT_22B_SZ 288

`define URAM288E5__INIT_22C    32'h00000239
`define URAM288E5__INIT_22C_SZ 288

`define URAM288E5__INIT_22D    32'h0000023a
`define URAM288E5__INIT_22D_SZ 288

`define URAM288E5__INIT_22E    32'h0000023b
`define URAM288E5__INIT_22E_SZ 288

`define URAM288E5__INIT_22F    32'h0000023c
`define URAM288E5__INIT_22F_SZ 288

`define URAM288E5__INIT_230    32'h0000023d
`define URAM288E5__INIT_230_SZ 288

`define URAM288E5__INIT_231    32'h0000023e
`define URAM288E5__INIT_231_SZ 288

`define URAM288E5__INIT_232    32'h0000023f
`define URAM288E5__INIT_232_SZ 288

`define URAM288E5__INIT_233    32'h00000240
`define URAM288E5__INIT_233_SZ 288

`define URAM288E5__INIT_234    32'h00000241
`define URAM288E5__INIT_234_SZ 288

`define URAM288E5__INIT_235    32'h00000242
`define URAM288E5__INIT_235_SZ 288

`define URAM288E5__INIT_236    32'h00000243
`define URAM288E5__INIT_236_SZ 288

`define URAM288E5__INIT_237    32'h00000244
`define URAM288E5__INIT_237_SZ 288

`define URAM288E5__INIT_238    32'h00000245
`define URAM288E5__INIT_238_SZ 288

`define URAM288E5__INIT_239    32'h00000246
`define URAM288E5__INIT_239_SZ 288

`define URAM288E5__INIT_23A    32'h00000247
`define URAM288E5__INIT_23A_SZ 288

`define URAM288E5__INIT_23B    32'h00000248
`define URAM288E5__INIT_23B_SZ 288

`define URAM288E5__INIT_23C    32'h00000249
`define URAM288E5__INIT_23C_SZ 288

`define URAM288E5__INIT_23D    32'h0000024a
`define URAM288E5__INIT_23D_SZ 288

`define URAM288E5__INIT_23E    32'h0000024b
`define URAM288E5__INIT_23E_SZ 288

`define URAM288E5__INIT_23F    32'h0000024c
`define URAM288E5__INIT_23F_SZ 288

`define URAM288E5__INIT_240    32'h0000024d
`define URAM288E5__INIT_240_SZ 288

`define URAM288E5__INIT_241    32'h0000024e
`define URAM288E5__INIT_241_SZ 288

`define URAM288E5__INIT_242    32'h0000024f
`define URAM288E5__INIT_242_SZ 288

`define URAM288E5__INIT_243    32'h00000250
`define URAM288E5__INIT_243_SZ 288

`define URAM288E5__INIT_244    32'h00000251
`define URAM288E5__INIT_244_SZ 288

`define URAM288E5__INIT_245    32'h00000252
`define URAM288E5__INIT_245_SZ 288

`define URAM288E5__INIT_246    32'h00000253
`define URAM288E5__INIT_246_SZ 288

`define URAM288E5__INIT_247    32'h00000254
`define URAM288E5__INIT_247_SZ 288

`define URAM288E5__INIT_248    32'h00000255
`define URAM288E5__INIT_248_SZ 288

`define URAM288E5__INIT_249    32'h00000256
`define URAM288E5__INIT_249_SZ 288

`define URAM288E5__INIT_24A    32'h00000257
`define URAM288E5__INIT_24A_SZ 288

`define URAM288E5__INIT_24B    32'h00000258
`define URAM288E5__INIT_24B_SZ 288

`define URAM288E5__INIT_24C    32'h00000259
`define URAM288E5__INIT_24C_SZ 288

`define URAM288E5__INIT_24D    32'h0000025a
`define URAM288E5__INIT_24D_SZ 288

`define URAM288E5__INIT_24E    32'h0000025b
`define URAM288E5__INIT_24E_SZ 288

`define URAM288E5__INIT_24F    32'h0000025c
`define URAM288E5__INIT_24F_SZ 288

`define URAM288E5__INIT_250    32'h0000025d
`define URAM288E5__INIT_250_SZ 288

`define URAM288E5__INIT_251    32'h0000025e
`define URAM288E5__INIT_251_SZ 288

`define URAM288E5__INIT_252    32'h0000025f
`define URAM288E5__INIT_252_SZ 288

`define URAM288E5__INIT_253    32'h00000260
`define URAM288E5__INIT_253_SZ 288

`define URAM288E5__INIT_254    32'h00000261
`define URAM288E5__INIT_254_SZ 288

`define URAM288E5__INIT_255    32'h00000262
`define URAM288E5__INIT_255_SZ 288

`define URAM288E5__INIT_256    32'h00000263
`define URAM288E5__INIT_256_SZ 288

`define URAM288E5__INIT_257    32'h00000264
`define URAM288E5__INIT_257_SZ 288

`define URAM288E5__INIT_258    32'h00000265
`define URAM288E5__INIT_258_SZ 288

`define URAM288E5__INIT_259    32'h00000266
`define URAM288E5__INIT_259_SZ 288

`define URAM288E5__INIT_25A    32'h00000267
`define URAM288E5__INIT_25A_SZ 288

`define URAM288E5__INIT_25B    32'h00000268
`define URAM288E5__INIT_25B_SZ 288

`define URAM288E5__INIT_25C    32'h00000269
`define URAM288E5__INIT_25C_SZ 288

`define URAM288E5__INIT_25D    32'h0000026a
`define URAM288E5__INIT_25D_SZ 288

`define URAM288E5__INIT_25E    32'h0000026b
`define URAM288E5__INIT_25E_SZ 288

`define URAM288E5__INIT_25F    32'h0000026c
`define URAM288E5__INIT_25F_SZ 288

`define URAM288E5__INIT_260    32'h0000026d
`define URAM288E5__INIT_260_SZ 288

`define URAM288E5__INIT_261    32'h0000026e
`define URAM288E5__INIT_261_SZ 288

`define URAM288E5__INIT_262    32'h0000026f
`define URAM288E5__INIT_262_SZ 288

`define URAM288E5__INIT_263    32'h00000270
`define URAM288E5__INIT_263_SZ 288

`define URAM288E5__INIT_264    32'h00000271
`define URAM288E5__INIT_264_SZ 288

`define URAM288E5__INIT_265    32'h00000272
`define URAM288E5__INIT_265_SZ 288

`define URAM288E5__INIT_266    32'h00000273
`define URAM288E5__INIT_266_SZ 288

`define URAM288E5__INIT_267    32'h00000274
`define URAM288E5__INIT_267_SZ 288

`define URAM288E5__INIT_268    32'h00000275
`define URAM288E5__INIT_268_SZ 288

`define URAM288E5__INIT_269    32'h00000276
`define URAM288E5__INIT_269_SZ 288

`define URAM288E5__INIT_26A    32'h00000277
`define URAM288E5__INIT_26A_SZ 288

`define URAM288E5__INIT_26B    32'h00000278
`define URAM288E5__INIT_26B_SZ 288

`define URAM288E5__INIT_26C    32'h00000279
`define URAM288E5__INIT_26C_SZ 288

`define URAM288E5__INIT_26D    32'h0000027a
`define URAM288E5__INIT_26D_SZ 288

`define URAM288E5__INIT_26E    32'h0000027b
`define URAM288E5__INIT_26E_SZ 288

`define URAM288E5__INIT_26F    32'h0000027c
`define URAM288E5__INIT_26F_SZ 288

`define URAM288E5__INIT_270    32'h0000027d
`define URAM288E5__INIT_270_SZ 288

`define URAM288E5__INIT_271    32'h0000027e
`define URAM288E5__INIT_271_SZ 288

`define URAM288E5__INIT_272    32'h0000027f
`define URAM288E5__INIT_272_SZ 288

`define URAM288E5__INIT_273    32'h00000280
`define URAM288E5__INIT_273_SZ 288

`define URAM288E5__INIT_274    32'h00000281
`define URAM288E5__INIT_274_SZ 288

`define URAM288E5__INIT_275    32'h00000282
`define URAM288E5__INIT_275_SZ 288

`define URAM288E5__INIT_276    32'h00000283
`define URAM288E5__INIT_276_SZ 288

`define URAM288E5__INIT_277    32'h00000284
`define URAM288E5__INIT_277_SZ 288

`define URAM288E5__INIT_278    32'h00000285
`define URAM288E5__INIT_278_SZ 288

`define URAM288E5__INIT_279    32'h00000286
`define URAM288E5__INIT_279_SZ 288

`define URAM288E5__INIT_27A    32'h00000287
`define URAM288E5__INIT_27A_SZ 288

`define URAM288E5__INIT_27B    32'h00000288
`define URAM288E5__INIT_27B_SZ 288

`define URAM288E5__INIT_27C    32'h00000289
`define URAM288E5__INIT_27C_SZ 288

`define URAM288E5__INIT_27D    32'h0000028a
`define URAM288E5__INIT_27D_SZ 288

`define URAM288E5__INIT_27E    32'h0000028b
`define URAM288E5__INIT_27E_SZ 288

`define URAM288E5__INIT_27F    32'h0000028c
`define URAM288E5__INIT_27F_SZ 288

`define URAM288E5__INIT_280    32'h0000028d
`define URAM288E5__INIT_280_SZ 288

`define URAM288E5__INIT_281    32'h0000028e
`define URAM288E5__INIT_281_SZ 288

`define URAM288E5__INIT_282    32'h0000028f
`define URAM288E5__INIT_282_SZ 288

`define URAM288E5__INIT_283    32'h00000290
`define URAM288E5__INIT_283_SZ 288

`define URAM288E5__INIT_284    32'h00000291
`define URAM288E5__INIT_284_SZ 288

`define URAM288E5__INIT_285    32'h00000292
`define URAM288E5__INIT_285_SZ 288

`define URAM288E5__INIT_286    32'h00000293
`define URAM288E5__INIT_286_SZ 288

`define URAM288E5__INIT_287    32'h00000294
`define URAM288E5__INIT_287_SZ 288

`define URAM288E5__INIT_288    32'h00000295
`define URAM288E5__INIT_288_SZ 288

`define URAM288E5__INIT_289    32'h00000296
`define URAM288E5__INIT_289_SZ 288

`define URAM288E5__INIT_28A    32'h00000297
`define URAM288E5__INIT_28A_SZ 288

`define URAM288E5__INIT_28B    32'h00000298
`define URAM288E5__INIT_28B_SZ 288

`define URAM288E5__INIT_28C    32'h00000299
`define URAM288E5__INIT_28C_SZ 288

`define URAM288E5__INIT_28D    32'h0000029a
`define URAM288E5__INIT_28D_SZ 288

`define URAM288E5__INIT_28E    32'h0000029b
`define URAM288E5__INIT_28E_SZ 288

`define URAM288E5__INIT_28F    32'h0000029c
`define URAM288E5__INIT_28F_SZ 288

`define URAM288E5__INIT_290    32'h0000029d
`define URAM288E5__INIT_290_SZ 288

`define URAM288E5__INIT_291    32'h0000029e
`define URAM288E5__INIT_291_SZ 288

`define URAM288E5__INIT_292    32'h0000029f
`define URAM288E5__INIT_292_SZ 288

`define URAM288E5__INIT_293    32'h000002a0
`define URAM288E5__INIT_293_SZ 288

`define URAM288E5__INIT_294    32'h000002a1
`define URAM288E5__INIT_294_SZ 288

`define URAM288E5__INIT_295    32'h000002a2
`define URAM288E5__INIT_295_SZ 288

`define URAM288E5__INIT_296    32'h000002a3
`define URAM288E5__INIT_296_SZ 288

`define URAM288E5__INIT_297    32'h000002a4
`define URAM288E5__INIT_297_SZ 288

`define URAM288E5__INIT_298    32'h000002a5
`define URAM288E5__INIT_298_SZ 288

`define URAM288E5__INIT_299    32'h000002a6
`define URAM288E5__INIT_299_SZ 288

`define URAM288E5__INIT_29A    32'h000002a7
`define URAM288E5__INIT_29A_SZ 288

`define URAM288E5__INIT_29B    32'h000002a8
`define URAM288E5__INIT_29B_SZ 288

`define URAM288E5__INIT_29C    32'h000002a9
`define URAM288E5__INIT_29C_SZ 288

`define URAM288E5__INIT_29D    32'h000002aa
`define URAM288E5__INIT_29D_SZ 288

`define URAM288E5__INIT_29E    32'h000002ab
`define URAM288E5__INIT_29E_SZ 288

`define URAM288E5__INIT_29F    32'h000002ac
`define URAM288E5__INIT_29F_SZ 288

`define URAM288E5__INIT_2A0    32'h000002ad
`define URAM288E5__INIT_2A0_SZ 288

`define URAM288E5__INIT_2A1    32'h000002ae
`define URAM288E5__INIT_2A1_SZ 288

`define URAM288E5__INIT_2A2    32'h000002af
`define URAM288E5__INIT_2A2_SZ 288

`define URAM288E5__INIT_2A3    32'h000002b0
`define URAM288E5__INIT_2A3_SZ 288

`define URAM288E5__INIT_2A4    32'h000002b1
`define URAM288E5__INIT_2A4_SZ 288

`define URAM288E5__INIT_2A5    32'h000002b2
`define URAM288E5__INIT_2A5_SZ 288

`define URAM288E5__INIT_2A6    32'h000002b3
`define URAM288E5__INIT_2A6_SZ 288

`define URAM288E5__INIT_2A7    32'h000002b4
`define URAM288E5__INIT_2A7_SZ 288

`define URAM288E5__INIT_2A8    32'h000002b5
`define URAM288E5__INIT_2A8_SZ 288

`define URAM288E5__INIT_2A9    32'h000002b6
`define URAM288E5__INIT_2A9_SZ 288

`define URAM288E5__INIT_2AA    32'h000002b7
`define URAM288E5__INIT_2AA_SZ 288

`define URAM288E5__INIT_2AB    32'h000002b8
`define URAM288E5__INIT_2AB_SZ 288

`define URAM288E5__INIT_2AC    32'h000002b9
`define URAM288E5__INIT_2AC_SZ 288

`define URAM288E5__INIT_2AD    32'h000002ba
`define URAM288E5__INIT_2AD_SZ 288

`define URAM288E5__INIT_2AE    32'h000002bb
`define URAM288E5__INIT_2AE_SZ 288

`define URAM288E5__INIT_2AF    32'h000002bc
`define URAM288E5__INIT_2AF_SZ 288

`define URAM288E5__INIT_2B0    32'h000002bd
`define URAM288E5__INIT_2B0_SZ 288

`define URAM288E5__INIT_2B1    32'h000002be
`define URAM288E5__INIT_2B1_SZ 288

`define URAM288E5__INIT_2B2    32'h000002bf
`define URAM288E5__INIT_2B2_SZ 288

`define URAM288E5__INIT_2B3    32'h000002c0
`define URAM288E5__INIT_2B3_SZ 288

`define URAM288E5__INIT_2B4    32'h000002c1
`define URAM288E5__INIT_2B4_SZ 288

`define URAM288E5__INIT_2B5    32'h000002c2
`define URAM288E5__INIT_2B5_SZ 288

`define URAM288E5__INIT_2B6    32'h000002c3
`define URAM288E5__INIT_2B6_SZ 288

`define URAM288E5__INIT_2B7    32'h000002c4
`define URAM288E5__INIT_2B7_SZ 288

`define URAM288E5__INIT_2B8    32'h000002c5
`define URAM288E5__INIT_2B8_SZ 288

`define URAM288E5__INIT_2B9    32'h000002c6
`define URAM288E5__INIT_2B9_SZ 288

`define URAM288E5__INIT_2BA    32'h000002c7
`define URAM288E5__INIT_2BA_SZ 288

`define URAM288E5__INIT_2BB    32'h000002c8
`define URAM288E5__INIT_2BB_SZ 288

`define URAM288E5__INIT_2BC    32'h000002c9
`define URAM288E5__INIT_2BC_SZ 288

`define URAM288E5__INIT_2BD    32'h000002ca
`define URAM288E5__INIT_2BD_SZ 288

`define URAM288E5__INIT_2BE    32'h000002cb
`define URAM288E5__INIT_2BE_SZ 288

`define URAM288E5__INIT_2BF    32'h000002cc
`define URAM288E5__INIT_2BF_SZ 288

`define URAM288E5__INIT_2C0    32'h000002cd
`define URAM288E5__INIT_2C0_SZ 288

`define URAM288E5__INIT_2C1    32'h000002ce
`define URAM288E5__INIT_2C1_SZ 288

`define URAM288E5__INIT_2C2    32'h000002cf
`define URAM288E5__INIT_2C2_SZ 288

`define URAM288E5__INIT_2C3    32'h000002d0
`define URAM288E5__INIT_2C3_SZ 288

`define URAM288E5__INIT_2C4    32'h000002d1
`define URAM288E5__INIT_2C4_SZ 288

`define URAM288E5__INIT_2C5    32'h000002d2
`define URAM288E5__INIT_2C5_SZ 288

`define URAM288E5__INIT_2C6    32'h000002d3
`define URAM288E5__INIT_2C6_SZ 288

`define URAM288E5__INIT_2C7    32'h000002d4
`define URAM288E5__INIT_2C7_SZ 288

`define URAM288E5__INIT_2C8    32'h000002d5
`define URAM288E5__INIT_2C8_SZ 288

`define URAM288E5__INIT_2C9    32'h000002d6
`define URAM288E5__INIT_2C9_SZ 288

`define URAM288E5__INIT_2CA    32'h000002d7
`define URAM288E5__INIT_2CA_SZ 288

`define URAM288E5__INIT_2CB    32'h000002d8
`define URAM288E5__INIT_2CB_SZ 288

`define URAM288E5__INIT_2CC    32'h000002d9
`define URAM288E5__INIT_2CC_SZ 288

`define URAM288E5__INIT_2CD    32'h000002da
`define URAM288E5__INIT_2CD_SZ 288

`define URAM288E5__INIT_2CE    32'h000002db
`define URAM288E5__INIT_2CE_SZ 288

`define URAM288E5__INIT_2CF    32'h000002dc
`define URAM288E5__INIT_2CF_SZ 288

`define URAM288E5__INIT_2D0    32'h000002dd
`define URAM288E5__INIT_2D0_SZ 288

`define URAM288E5__INIT_2D1    32'h000002de
`define URAM288E5__INIT_2D1_SZ 288

`define URAM288E5__INIT_2D2    32'h000002df
`define URAM288E5__INIT_2D2_SZ 288

`define URAM288E5__INIT_2D3    32'h000002e0
`define URAM288E5__INIT_2D3_SZ 288

`define URAM288E5__INIT_2D4    32'h000002e1
`define URAM288E5__INIT_2D4_SZ 288

`define URAM288E5__INIT_2D5    32'h000002e2
`define URAM288E5__INIT_2D5_SZ 288

`define URAM288E5__INIT_2D6    32'h000002e3
`define URAM288E5__INIT_2D6_SZ 288

`define URAM288E5__INIT_2D7    32'h000002e4
`define URAM288E5__INIT_2D7_SZ 288

`define URAM288E5__INIT_2D8    32'h000002e5
`define URAM288E5__INIT_2D8_SZ 288

`define URAM288E5__INIT_2D9    32'h000002e6
`define URAM288E5__INIT_2D9_SZ 288

`define URAM288E5__INIT_2DA    32'h000002e7
`define URAM288E5__INIT_2DA_SZ 288

`define URAM288E5__INIT_2DB    32'h000002e8
`define URAM288E5__INIT_2DB_SZ 288

`define URAM288E5__INIT_2DC    32'h000002e9
`define URAM288E5__INIT_2DC_SZ 288

`define URAM288E5__INIT_2DD    32'h000002ea
`define URAM288E5__INIT_2DD_SZ 288

`define URAM288E5__INIT_2DE    32'h000002eb
`define URAM288E5__INIT_2DE_SZ 288

`define URAM288E5__INIT_2DF    32'h000002ec
`define URAM288E5__INIT_2DF_SZ 288

`define URAM288E5__INIT_2E0    32'h000002ed
`define URAM288E5__INIT_2E0_SZ 288

`define URAM288E5__INIT_2E1    32'h000002ee
`define URAM288E5__INIT_2E1_SZ 288

`define URAM288E5__INIT_2E2    32'h000002ef
`define URAM288E5__INIT_2E2_SZ 288

`define URAM288E5__INIT_2E3    32'h000002f0
`define URAM288E5__INIT_2E3_SZ 288

`define URAM288E5__INIT_2E4    32'h000002f1
`define URAM288E5__INIT_2E4_SZ 288

`define URAM288E5__INIT_2E5    32'h000002f2
`define URAM288E5__INIT_2E5_SZ 288

`define URAM288E5__INIT_2E6    32'h000002f3
`define URAM288E5__INIT_2E6_SZ 288

`define URAM288E5__INIT_2E7    32'h000002f4
`define URAM288E5__INIT_2E7_SZ 288

`define URAM288E5__INIT_2E8    32'h000002f5
`define URAM288E5__INIT_2E8_SZ 288

`define URAM288E5__INIT_2E9    32'h000002f6
`define URAM288E5__INIT_2E9_SZ 288

`define URAM288E5__INIT_2EA    32'h000002f7
`define URAM288E5__INIT_2EA_SZ 288

`define URAM288E5__INIT_2EB    32'h000002f8
`define URAM288E5__INIT_2EB_SZ 288

`define URAM288E5__INIT_2EC    32'h000002f9
`define URAM288E5__INIT_2EC_SZ 288

`define URAM288E5__INIT_2ED    32'h000002fa
`define URAM288E5__INIT_2ED_SZ 288

`define URAM288E5__INIT_2EE    32'h000002fb
`define URAM288E5__INIT_2EE_SZ 288

`define URAM288E5__INIT_2EF    32'h000002fc
`define URAM288E5__INIT_2EF_SZ 288

`define URAM288E5__INIT_2F0    32'h000002fd
`define URAM288E5__INIT_2F0_SZ 288

`define URAM288E5__INIT_2F1    32'h000002fe
`define URAM288E5__INIT_2F1_SZ 288

`define URAM288E5__INIT_2F2    32'h000002ff
`define URAM288E5__INIT_2F2_SZ 288

`define URAM288E5__INIT_2F3    32'h00000300
`define URAM288E5__INIT_2F3_SZ 288

`define URAM288E5__INIT_2F4    32'h00000301
`define URAM288E5__INIT_2F4_SZ 288

`define URAM288E5__INIT_2F5    32'h00000302
`define URAM288E5__INIT_2F5_SZ 288

`define URAM288E5__INIT_2F6    32'h00000303
`define URAM288E5__INIT_2F6_SZ 288

`define URAM288E5__INIT_2F7    32'h00000304
`define URAM288E5__INIT_2F7_SZ 288

`define URAM288E5__INIT_2F8    32'h00000305
`define URAM288E5__INIT_2F8_SZ 288

`define URAM288E5__INIT_2F9    32'h00000306
`define URAM288E5__INIT_2F9_SZ 288

`define URAM288E5__INIT_2FA    32'h00000307
`define URAM288E5__INIT_2FA_SZ 288

`define URAM288E5__INIT_2FB    32'h00000308
`define URAM288E5__INIT_2FB_SZ 288

`define URAM288E5__INIT_2FC    32'h00000309
`define URAM288E5__INIT_2FC_SZ 288

`define URAM288E5__INIT_2FD    32'h0000030a
`define URAM288E5__INIT_2FD_SZ 288

`define URAM288E5__INIT_2FE    32'h0000030b
`define URAM288E5__INIT_2FE_SZ 288

`define URAM288E5__INIT_2FF    32'h0000030c
`define URAM288E5__INIT_2FF_SZ 288

`define URAM288E5__INIT_300    32'h0000030d
`define URAM288E5__INIT_300_SZ 288

`define URAM288E5__INIT_301    32'h0000030e
`define URAM288E5__INIT_301_SZ 288

`define URAM288E5__INIT_302    32'h0000030f
`define URAM288E5__INIT_302_SZ 288

`define URAM288E5__INIT_303    32'h00000310
`define URAM288E5__INIT_303_SZ 288

`define URAM288E5__INIT_304    32'h00000311
`define URAM288E5__INIT_304_SZ 288

`define URAM288E5__INIT_305    32'h00000312
`define URAM288E5__INIT_305_SZ 288

`define URAM288E5__INIT_306    32'h00000313
`define URAM288E5__INIT_306_SZ 288

`define URAM288E5__INIT_307    32'h00000314
`define URAM288E5__INIT_307_SZ 288

`define URAM288E5__INIT_308    32'h00000315
`define URAM288E5__INIT_308_SZ 288

`define URAM288E5__INIT_309    32'h00000316
`define URAM288E5__INIT_309_SZ 288

`define URAM288E5__INIT_30A    32'h00000317
`define URAM288E5__INIT_30A_SZ 288

`define URAM288E5__INIT_30B    32'h00000318
`define URAM288E5__INIT_30B_SZ 288

`define URAM288E5__INIT_30C    32'h00000319
`define URAM288E5__INIT_30C_SZ 288

`define URAM288E5__INIT_30D    32'h0000031a
`define URAM288E5__INIT_30D_SZ 288

`define URAM288E5__INIT_30E    32'h0000031b
`define URAM288E5__INIT_30E_SZ 288

`define URAM288E5__INIT_30F    32'h0000031c
`define URAM288E5__INIT_30F_SZ 288

`define URAM288E5__INIT_310    32'h0000031d
`define URAM288E5__INIT_310_SZ 288

`define URAM288E5__INIT_311    32'h0000031e
`define URAM288E5__INIT_311_SZ 288

`define URAM288E5__INIT_312    32'h0000031f
`define URAM288E5__INIT_312_SZ 288

`define URAM288E5__INIT_313    32'h00000320
`define URAM288E5__INIT_313_SZ 288

`define URAM288E5__INIT_314    32'h00000321
`define URAM288E5__INIT_314_SZ 288

`define URAM288E5__INIT_315    32'h00000322
`define URAM288E5__INIT_315_SZ 288

`define URAM288E5__INIT_316    32'h00000323
`define URAM288E5__INIT_316_SZ 288

`define URAM288E5__INIT_317    32'h00000324
`define URAM288E5__INIT_317_SZ 288

`define URAM288E5__INIT_318    32'h00000325
`define URAM288E5__INIT_318_SZ 288

`define URAM288E5__INIT_319    32'h00000326
`define URAM288E5__INIT_319_SZ 288

`define URAM288E5__INIT_31A    32'h00000327
`define URAM288E5__INIT_31A_SZ 288

`define URAM288E5__INIT_31B    32'h00000328
`define URAM288E5__INIT_31B_SZ 288

`define URAM288E5__INIT_31C    32'h00000329
`define URAM288E5__INIT_31C_SZ 288

`define URAM288E5__INIT_31D    32'h0000032a
`define URAM288E5__INIT_31D_SZ 288

`define URAM288E5__INIT_31E    32'h0000032b
`define URAM288E5__INIT_31E_SZ 288

`define URAM288E5__INIT_31F    32'h0000032c
`define URAM288E5__INIT_31F_SZ 288

`define URAM288E5__INIT_320    32'h0000032d
`define URAM288E5__INIT_320_SZ 288

`define URAM288E5__INIT_321    32'h0000032e
`define URAM288E5__INIT_321_SZ 288

`define URAM288E5__INIT_322    32'h0000032f
`define URAM288E5__INIT_322_SZ 288

`define URAM288E5__INIT_323    32'h00000330
`define URAM288E5__INIT_323_SZ 288

`define URAM288E5__INIT_324    32'h00000331
`define URAM288E5__INIT_324_SZ 288

`define URAM288E5__INIT_325    32'h00000332
`define URAM288E5__INIT_325_SZ 288

`define URAM288E5__INIT_326    32'h00000333
`define URAM288E5__INIT_326_SZ 288

`define URAM288E5__INIT_327    32'h00000334
`define URAM288E5__INIT_327_SZ 288

`define URAM288E5__INIT_328    32'h00000335
`define URAM288E5__INIT_328_SZ 288

`define URAM288E5__INIT_329    32'h00000336
`define URAM288E5__INIT_329_SZ 288

`define URAM288E5__INIT_32A    32'h00000337
`define URAM288E5__INIT_32A_SZ 288

`define URAM288E5__INIT_32B    32'h00000338
`define URAM288E5__INIT_32B_SZ 288

`define URAM288E5__INIT_32C    32'h00000339
`define URAM288E5__INIT_32C_SZ 288

`define URAM288E5__INIT_32D    32'h0000033a
`define URAM288E5__INIT_32D_SZ 288

`define URAM288E5__INIT_32E    32'h0000033b
`define URAM288E5__INIT_32E_SZ 288

`define URAM288E5__INIT_32F    32'h0000033c
`define URAM288E5__INIT_32F_SZ 288

`define URAM288E5__INIT_330    32'h0000033d
`define URAM288E5__INIT_330_SZ 288

`define URAM288E5__INIT_331    32'h0000033e
`define URAM288E5__INIT_331_SZ 288

`define URAM288E5__INIT_332    32'h0000033f
`define URAM288E5__INIT_332_SZ 288

`define URAM288E5__INIT_333    32'h00000340
`define URAM288E5__INIT_333_SZ 288

`define URAM288E5__INIT_334    32'h00000341
`define URAM288E5__INIT_334_SZ 288

`define URAM288E5__INIT_335    32'h00000342
`define URAM288E5__INIT_335_SZ 288

`define URAM288E5__INIT_336    32'h00000343
`define URAM288E5__INIT_336_SZ 288

`define URAM288E5__INIT_337    32'h00000344
`define URAM288E5__INIT_337_SZ 288

`define URAM288E5__INIT_338    32'h00000345
`define URAM288E5__INIT_338_SZ 288

`define URAM288E5__INIT_339    32'h00000346
`define URAM288E5__INIT_339_SZ 288

`define URAM288E5__INIT_33A    32'h00000347
`define URAM288E5__INIT_33A_SZ 288

`define URAM288E5__INIT_33B    32'h00000348
`define URAM288E5__INIT_33B_SZ 288

`define URAM288E5__INIT_33C    32'h00000349
`define URAM288E5__INIT_33C_SZ 288

`define URAM288E5__INIT_33D    32'h0000034a
`define URAM288E5__INIT_33D_SZ 288

`define URAM288E5__INIT_33E    32'h0000034b
`define URAM288E5__INIT_33E_SZ 288

`define URAM288E5__INIT_33F    32'h0000034c
`define URAM288E5__INIT_33F_SZ 288

`define URAM288E5__INIT_340    32'h0000034d
`define URAM288E5__INIT_340_SZ 288

`define URAM288E5__INIT_341    32'h0000034e
`define URAM288E5__INIT_341_SZ 288

`define URAM288E5__INIT_342    32'h0000034f
`define URAM288E5__INIT_342_SZ 288

`define URAM288E5__INIT_343    32'h00000350
`define URAM288E5__INIT_343_SZ 288

`define URAM288E5__INIT_344    32'h00000351
`define URAM288E5__INIT_344_SZ 288

`define URAM288E5__INIT_345    32'h00000352
`define URAM288E5__INIT_345_SZ 288

`define URAM288E5__INIT_346    32'h00000353
`define URAM288E5__INIT_346_SZ 288

`define URAM288E5__INIT_347    32'h00000354
`define URAM288E5__INIT_347_SZ 288

`define URAM288E5__INIT_348    32'h00000355
`define URAM288E5__INIT_348_SZ 288

`define URAM288E5__INIT_349    32'h00000356
`define URAM288E5__INIT_349_SZ 288

`define URAM288E5__INIT_34A    32'h00000357
`define URAM288E5__INIT_34A_SZ 288

`define URAM288E5__INIT_34B    32'h00000358
`define URAM288E5__INIT_34B_SZ 288

`define URAM288E5__INIT_34C    32'h00000359
`define URAM288E5__INIT_34C_SZ 288

`define URAM288E5__INIT_34D    32'h0000035a
`define URAM288E5__INIT_34D_SZ 288

`define URAM288E5__INIT_34E    32'h0000035b
`define URAM288E5__INIT_34E_SZ 288

`define URAM288E5__INIT_34F    32'h0000035c
`define URAM288E5__INIT_34F_SZ 288

`define URAM288E5__INIT_350    32'h0000035d
`define URAM288E5__INIT_350_SZ 288

`define URAM288E5__INIT_351    32'h0000035e
`define URAM288E5__INIT_351_SZ 288

`define URAM288E5__INIT_352    32'h0000035f
`define URAM288E5__INIT_352_SZ 288

`define URAM288E5__INIT_353    32'h00000360
`define URAM288E5__INIT_353_SZ 288

`define URAM288E5__INIT_354    32'h00000361
`define URAM288E5__INIT_354_SZ 288

`define URAM288E5__INIT_355    32'h00000362
`define URAM288E5__INIT_355_SZ 288

`define URAM288E5__INIT_356    32'h00000363
`define URAM288E5__INIT_356_SZ 288

`define URAM288E5__INIT_357    32'h00000364
`define URAM288E5__INIT_357_SZ 288

`define URAM288E5__INIT_358    32'h00000365
`define URAM288E5__INIT_358_SZ 288

`define URAM288E5__INIT_359    32'h00000366
`define URAM288E5__INIT_359_SZ 288

`define URAM288E5__INIT_35A    32'h00000367
`define URAM288E5__INIT_35A_SZ 288

`define URAM288E5__INIT_35B    32'h00000368
`define URAM288E5__INIT_35B_SZ 288

`define URAM288E5__INIT_35C    32'h00000369
`define URAM288E5__INIT_35C_SZ 288

`define URAM288E5__INIT_35D    32'h0000036a
`define URAM288E5__INIT_35D_SZ 288

`define URAM288E5__INIT_35E    32'h0000036b
`define URAM288E5__INIT_35E_SZ 288

`define URAM288E5__INIT_35F    32'h0000036c
`define URAM288E5__INIT_35F_SZ 288

`define URAM288E5__INIT_360    32'h0000036d
`define URAM288E5__INIT_360_SZ 288

`define URAM288E5__INIT_361    32'h0000036e
`define URAM288E5__INIT_361_SZ 288

`define URAM288E5__INIT_362    32'h0000036f
`define URAM288E5__INIT_362_SZ 288

`define URAM288E5__INIT_363    32'h00000370
`define URAM288E5__INIT_363_SZ 288

`define URAM288E5__INIT_364    32'h00000371
`define URAM288E5__INIT_364_SZ 288

`define URAM288E5__INIT_365    32'h00000372
`define URAM288E5__INIT_365_SZ 288

`define URAM288E5__INIT_366    32'h00000373
`define URAM288E5__INIT_366_SZ 288

`define URAM288E5__INIT_367    32'h00000374
`define URAM288E5__INIT_367_SZ 288

`define URAM288E5__INIT_368    32'h00000375
`define URAM288E5__INIT_368_SZ 288

`define URAM288E5__INIT_369    32'h00000376
`define URAM288E5__INIT_369_SZ 288

`define URAM288E5__INIT_36A    32'h00000377
`define URAM288E5__INIT_36A_SZ 288

`define URAM288E5__INIT_36B    32'h00000378
`define URAM288E5__INIT_36B_SZ 288

`define URAM288E5__INIT_36C    32'h00000379
`define URAM288E5__INIT_36C_SZ 288

`define URAM288E5__INIT_36D    32'h0000037a
`define URAM288E5__INIT_36D_SZ 288

`define URAM288E5__INIT_36E    32'h0000037b
`define URAM288E5__INIT_36E_SZ 288

`define URAM288E5__INIT_36F    32'h0000037c
`define URAM288E5__INIT_36F_SZ 288

`define URAM288E5__INIT_370    32'h0000037d
`define URAM288E5__INIT_370_SZ 288

`define URAM288E5__INIT_371    32'h0000037e
`define URAM288E5__INIT_371_SZ 288

`define URAM288E5__INIT_372    32'h0000037f
`define URAM288E5__INIT_372_SZ 288

`define URAM288E5__INIT_373    32'h00000380
`define URAM288E5__INIT_373_SZ 288

`define URAM288E5__INIT_374    32'h00000381
`define URAM288E5__INIT_374_SZ 288

`define URAM288E5__INIT_375    32'h00000382
`define URAM288E5__INIT_375_SZ 288

`define URAM288E5__INIT_376    32'h00000383
`define URAM288E5__INIT_376_SZ 288

`define URAM288E5__INIT_377    32'h00000384
`define URAM288E5__INIT_377_SZ 288

`define URAM288E5__INIT_378    32'h00000385
`define URAM288E5__INIT_378_SZ 288

`define URAM288E5__INIT_379    32'h00000386
`define URAM288E5__INIT_379_SZ 288

`define URAM288E5__INIT_37A    32'h00000387
`define URAM288E5__INIT_37A_SZ 288

`define URAM288E5__INIT_37B    32'h00000388
`define URAM288E5__INIT_37B_SZ 288

`define URAM288E5__INIT_37C    32'h00000389
`define URAM288E5__INIT_37C_SZ 288

`define URAM288E5__INIT_37D    32'h0000038a
`define URAM288E5__INIT_37D_SZ 288

`define URAM288E5__INIT_37E    32'h0000038b
`define URAM288E5__INIT_37E_SZ 288

`define URAM288E5__INIT_37F    32'h0000038c
`define URAM288E5__INIT_37F_SZ 288

`define URAM288E5__INIT_380    32'h0000038d
`define URAM288E5__INIT_380_SZ 288

`define URAM288E5__INIT_381    32'h0000038e
`define URAM288E5__INIT_381_SZ 288

`define URAM288E5__INIT_382    32'h0000038f
`define URAM288E5__INIT_382_SZ 288

`define URAM288E5__INIT_383    32'h00000390
`define URAM288E5__INIT_383_SZ 288

`define URAM288E5__INIT_384    32'h00000391
`define URAM288E5__INIT_384_SZ 288

`define URAM288E5__INIT_385    32'h00000392
`define URAM288E5__INIT_385_SZ 288

`define URAM288E5__INIT_386    32'h00000393
`define URAM288E5__INIT_386_SZ 288

`define URAM288E5__INIT_387    32'h00000394
`define URAM288E5__INIT_387_SZ 288

`define URAM288E5__INIT_388    32'h00000395
`define URAM288E5__INIT_388_SZ 288

`define URAM288E5__INIT_389    32'h00000396
`define URAM288E5__INIT_389_SZ 288

`define URAM288E5__INIT_38A    32'h00000397
`define URAM288E5__INIT_38A_SZ 288

`define URAM288E5__INIT_38B    32'h00000398
`define URAM288E5__INIT_38B_SZ 288

`define URAM288E5__INIT_38C    32'h00000399
`define URAM288E5__INIT_38C_SZ 288

`define URAM288E5__INIT_38D    32'h0000039a
`define URAM288E5__INIT_38D_SZ 288

`define URAM288E5__INIT_38E    32'h0000039b
`define URAM288E5__INIT_38E_SZ 288

`define URAM288E5__INIT_38F    32'h0000039c
`define URAM288E5__INIT_38F_SZ 288

`define URAM288E5__INIT_390    32'h0000039d
`define URAM288E5__INIT_390_SZ 288

`define URAM288E5__INIT_391    32'h0000039e
`define URAM288E5__INIT_391_SZ 288

`define URAM288E5__INIT_392    32'h0000039f
`define URAM288E5__INIT_392_SZ 288

`define URAM288E5__INIT_393    32'h000003a0
`define URAM288E5__INIT_393_SZ 288

`define URAM288E5__INIT_394    32'h000003a1
`define URAM288E5__INIT_394_SZ 288

`define URAM288E5__INIT_395    32'h000003a2
`define URAM288E5__INIT_395_SZ 288

`define URAM288E5__INIT_396    32'h000003a3
`define URAM288E5__INIT_396_SZ 288

`define URAM288E5__INIT_397    32'h000003a4
`define URAM288E5__INIT_397_SZ 288

`define URAM288E5__INIT_398    32'h000003a5
`define URAM288E5__INIT_398_SZ 288

`define URAM288E5__INIT_399    32'h000003a6
`define URAM288E5__INIT_399_SZ 288

`define URAM288E5__INIT_39A    32'h000003a7
`define URAM288E5__INIT_39A_SZ 288

`define URAM288E5__INIT_39B    32'h000003a8
`define URAM288E5__INIT_39B_SZ 288

`define URAM288E5__INIT_39C    32'h000003a9
`define URAM288E5__INIT_39C_SZ 288

`define URAM288E5__INIT_39D    32'h000003aa
`define URAM288E5__INIT_39D_SZ 288

`define URAM288E5__INIT_39E    32'h000003ab
`define URAM288E5__INIT_39E_SZ 288

`define URAM288E5__INIT_39F    32'h000003ac
`define URAM288E5__INIT_39F_SZ 288

`define URAM288E5__INIT_3A0    32'h000003ad
`define URAM288E5__INIT_3A0_SZ 288

`define URAM288E5__INIT_3A1    32'h000003ae
`define URAM288E5__INIT_3A1_SZ 288

`define URAM288E5__INIT_3A2    32'h000003af
`define URAM288E5__INIT_3A2_SZ 288

`define URAM288E5__INIT_3A3    32'h000003b0
`define URAM288E5__INIT_3A3_SZ 288

`define URAM288E5__INIT_3A4    32'h000003b1
`define URAM288E5__INIT_3A4_SZ 288

`define URAM288E5__INIT_3A5    32'h000003b2
`define URAM288E5__INIT_3A5_SZ 288

`define URAM288E5__INIT_3A6    32'h000003b3
`define URAM288E5__INIT_3A6_SZ 288

`define URAM288E5__INIT_3A7    32'h000003b4
`define URAM288E5__INIT_3A7_SZ 288

`define URAM288E5__INIT_3A8    32'h000003b5
`define URAM288E5__INIT_3A8_SZ 288

`define URAM288E5__INIT_3A9    32'h000003b6
`define URAM288E5__INIT_3A9_SZ 288

`define URAM288E5__INIT_3AA    32'h000003b7
`define URAM288E5__INIT_3AA_SZ 288

`define URAM288E5__INIT_3AB    32'h000003b8
`define URAM288E5__INIT_3AB_SZ 288

`define URAM288E5__INIT_3AC    32'h000003b9
`define URAM288E5__INIT_3AC_SZ 288

`define URAM288E5__INIT_3AD    32'h000003ba
`define URAM288E5__INIT_3AD_SZ 288

`define URAM288E5__INIT_3AE    32'h000003bb
`define URAM288E5__INIT_3AE_SZ 288

`define URAM288E5__INIT_3AF    32'h000003bc
`define URAM288E5__INIT_3AF_SZ 288

`define URAM288E5__INIT_3B0    32'h000003bd
`define URAM288E5__INIT_3B0_SZ 288

`define URAM288E5__INIT_3B1    32'h000003be
`define URAM288E5__INIT_3B1_SZ 288

`define URAM288E5__INIT_3B2    32'h000003bf
`define URAM288E5__INIT_3B2_SZ 288

`define URAM288E5__INIT_3B3    32'h000003c0
`define URAM288E5__INIT_3B3_SZ 288

`define URAM288E5__INIT_3B4    32'h000003c1
`define URAM288E5__INIT_3B4_SZ 288

`define URAM288E5__INIT_3B5    32'h000003c2
`define URAM288E5__INIT_3B5_SZ 288

`define URAM288E5__INIT_3B6    32'h000003c3
`define URAM288E5__INIT_3B6_SZ 288

`define URAM288E5__INIT_3B7    32'h000003c4
`define URAM288E5__INIT_3B7_SZ 288

`define URAM288E5__INIT_3B8    32'h000003c5
`define URAM288E5__INIT_3B8_SZ 288

`define URAM288E5__INIT_3B9    32'h000003c6
`define URAM288E5__INIT_3B9_SZ 288

`define URAM288E5__INIT_3BA    32'h000003c7
`define URAM288E5__INIT_3BA_SZ 288

`define URAM288E5__INIT_3BB    32'h000003c8
`define URAM288E5__INIT_3BB_SZ 288

`define URAM288E5__INIT_3BC    32'h000003c9
`define URAM288E5__INIT_3BC_SZ 288

`define URAM288E5__INIT_3BD    32'h000003ca
`define URAM288E5__INIT_3BD_SZ 288

`define URAM288E5__INIT_3BE    32'h000003cb
`define URAM288E5__INIT_3BE_SZ 288

`define URAM288E5__INIT_3BF    32'h000003cc
`define URAM288E5__INIT_3BF_SZ 288

`define URAM288E5__INIT_3C0    32'h000003cd
`define URAM288E5__INIT_3C0_SZ 288

`define URAM288E5__INIT_3C1    32'h000003ce
`define URAM288E5__INIT_3C1_SZ 288

`define URAM288E5__INIT_3C2    32'h000003cf
`define URAM288E5__INIT_3C2_SZ 288

`define URAM288E5__INIT_3C3    32'h000003d0
`define URAM288E5__INIT_3C3_SZ 288

`define URAM288E5__INIT_3C4    32'h000003d1
`define URAM288E5__INIT_3C4_SZ 288

`define URAM288E5__INIT_3C5    32'h000003d2
`define URAM288E5__INIT_3C5_SZ 288

`define URAM288E5__INIT_3C6    32'h000003d3
`define URAM288E5__INIT_3C6_SZ 288

`define URAM288E5__INIT_3C7    32'h000003d4
`define URAM288E5__INIT_3C7_SZ 288

`define URAM288E5__INIT_3C8    32'h000003d5
`define URAM288E5__INIT_3C8_SZ 288

`define URAM288E5__INIT_3C9    32'h000003d6
`define URAM288E5__INIT_3C9_SZ 288

`define URAM288E5__INIT_3CA    32'h000003d7
`define URAM288E5__INIT_3CA_SZ 288

`define URAM288E5__INIT_3CB    32'h000003d8
`define URAM288E5__INIT_3CB_SZ 288

`define URAM288E5__INIT_3CC    32'h000003d9
`define URAM288E5__INIT_3CC_SZ 288

`define URAM288E5__INIT_3CD    32'h000003da
`define URAM288E5__INIT_3CD_SZ 288

`define URAM288E5__INIT_3CE    32'h000003db
`define URAM288E5__INIT_3CE_SZ 288

`define URAM288E5__INIT_3CF    32'h000003dc
`define URAM288E5__INIT_3CF_SZ 288

`define URAM288E5__INIT_3D0    32'h000003dd
`define URAM288E5__INIT_3D0_SZ 288

`define URAM288E5__INIT_3D1    32'h000003de
`define URAM288E5__INIT_3D1_SZ 288

`define URAM288E5__INIT_3D2    32'h000003df
`define URAM288E5__INIT_3D2_SZ 288

`define URAM288E5__INIT_3D3    32'h000003e0
`define URAM288E5__INIT_3D3_SZ 288

`define URAM288E5__INIT_3D4    32'h000003e1
`define URAM288E5__INIT_3D4_SZ 288

`define URAM288E5__INIT_3D5    32'h000003e2
`define URAM288E5__INIT_3D5_SZ 288

`define URAM288E5__INIT_3D6    32'h000003e3
`define URAM288E5__INIT_3D6_SZ 288

`define URAM288E5__INIT_3D7    32'h000003e4
`define URAM288E5__INIT_3D7_SZ 288

`define URAM288E5__INIT_3D8    32'h000003e5
`define URAM288E5__INIT_3D8_SZ 288

`define URAM288E5__INIT_3D9    32'h000003e6
`define URAM288E5__INIT_3D9_SZ 288

`define URAM288E5__INIT_3DA    32'h000003e7
`define URAM288E5__INIT_3DA_SZ 288

`define URAM288E5__INIT_3DB    32'h000003e8
`define URAM288E5__INIT_3DB_SZ 288

`define URAM288E5__INIT_3DC    32'h000003e9
`define URAM288E5__INIT_3DC_SZ 288

`define URAM288E5__INIT_3DD    32'h000003ea
`define URAM288E5__INIT_3DD_SZ 288

`define URAM288E5__INIT_3DE    32'h000003eb
`define URAM288E5__INIT_3DE_SZ 288

`define URAM288E5__INIT_3DF    32'h000003ec
`define URAM288E5__INIT_3DF_SZ 288

`define URAM288E5__INIT_3E0    32'h000003ed
`define URAM288E5__INIT_3E0_SZ 288

`define URAM288E5__INIT_3E1    32'h000003ee
`define URAM288E5__INIT_3E1_SZ 288

`define URAM288E5__INIT_3E2    32'h000003ef
`define URAM288E5__INIT_3E2_SZ 288

`define URAM288E5__INIT_3E3    32'h000003f0
`define URAM288E5__INIT_3E3_SZ 288

`define URAM288E5__INIT_3E4    32'h000003f1
`define URAM288E5__INIT_3E4_SZ 288

`define URAM288E5__INIT_3E5    32'h000003f2
`define URAM288E5__INIT_3E5_SZ 288

`define URAM288E5__INIT_3E6    32'h000003f3
`define URAM288E5__INIT_3E6_SZ 288

`define URAM288E5__INIT_3E7    32'h000003f4
`define URAM288E5__INIT_3E7_SZ 288

`define URAM288E5__INIT_3E8    32'h000003f5
`define URAM288E5__INIT_3E8_SZ 288

`define URAM288E5__INIT_3E9    32'h000003f6
`define URAM288E5__INIT_3E9_SZ 288

`define URAM288E5__INIT_3EA    32'h000003f7
`define URAM288E5__INIT_3EA_SZ 288

`define URAM288E5__INIT_3EB    32'h000003f8
`define URAM288E5__INIT_3EB_SZ 288

`define URAM288E5__INIT_3EC    32'h000003f9
`define URAM288E5__INIT_3EC_SZ 288

`define URAM288E5__INIT_3ED    32'h000003fa
`define URAM288E5__INIT_3ED_SZ 288

`define URAM288E5__INIT_3EE    32'h000003fb
`define URAM288E5__INIT_3EE_SZ 288

`define URAM288E5__INIT_3EF    32'h000003fc
`define URAM288E5__INIT_3EF_SZ 288

`define URAM288E5__INIT_3F0    32'h000003fd
`define URAM288E5__INIT_3F0_SZ 288

`define URAM288E5__INIT_3F1    32'h000003fe
`define URAM288E5__INIT_3F1_SZ 288

`define URAM288E5__INIT_3F2    32'h000003ff
`define URAM288E5__INIT_3F2_SZ 288

`define URAM288E5__INIT_3F3    32'h00000400
`define URAM288E5__INIT_3F3_SZ 288

`define URAM288E5__INIT_3F4    32'h00000401
`define URAM288E5__INIT_3F4_SZ 288

`define URAM288E5__INIT_3F5    32'h00000402
`define URAM288E5__INIT_3F5_SZ 288

`define URAM288E5__INIT_3F6    32'h00000403
`define URAM288E5__INIT_3F6_SZ 288

`define URAM288E5__INIT_3F7    32'h00000404
`define URAM288E5__INIT_3F7_SZ 288

`define URAM288E5__INIT_3F8    32'h00000405
`define URAM288E5__INIT_3F8_SZ 288

`define URAM288E5__INIT_3F9    32'h00000406
`define URAM288E5__INIT_3F9_SZ 288

`define URAM288E5__INIT_3FA    32'h00000407
`define URAM288E5__INIT_3FA_SZ 288

`define URAM288E5__INIT_3FB    32'h00000408
`define URAM288E5__INIT_3FB_SZ 288

`define URAM288E5__INIT_3FC    32'h00000409
`define URAM288E5__INIT_3FC_SZ 288

`define URAM288E5__INIT_3FD    32'h0000040a
`define URAM288E5__INIT_3FD_SZ 288

`define URAM288E5__INIT_3FE    32'h0000040b
`define URAM288E5__INIT_3FE_SZ 288

`define URAM288E5__INIT_3FF    32'h0000040c
`define URAM288E5__INIT_3FF_SZ 288

`define URAM288E5__INIT_FILE    32'h0000040d
`define URAM288E5__INIT_FILE_SZ 32

`define URAM288E5__IREG_PRE_A    32'h0000040e
`define URAM288E5__IREG_PRE_A_SZ 40

`define URAM288E5__IREG_PRE_B    32'h0000040f
`define URAM288E5__IREG_PRE_B_SZ 40

`define URAM288E5__IS_CLK_INVERTED    32'h00000410
`define URAM288E5__IS_CLK_INVERTED_SZ 1

`define URAM288E5__IS_EN_A_INVERTED    32'h00000411
`define URAM288E5__IS_EN_A_INVERTED_SZ 1

`define URAM288E5__IS_EN_B_INVERTED    32'h00000412
`define URAM288E5__IS_EN_B_INVERTED_SZ 1

`define URAM288E5__IS_RDB_WR_A_INVERTED    32'h00000413
`define URAM288E5__IS_RDB_WR_A_INVERTED_SZ 1

`define URAM288E5__IS_RDB_WR_B_INVERTED    32'h00000414
`define URAM288E5__IS_RDB_WR_B_INVERTED_SZ 1

`define URAM288E5__IS_RST_A_INVERTED    32'h00000415
`define URAM288E5__IS_RST_A_INVERTED_SZ 1

`define URAM288E5__IS_RST_B_INVERTED    32'h00000416
`define URAM288E5__IS_RST_B_INVERTED_SZ 1

`define URAM288E5__MATRIX_ID    32'h00000417
`define URAM288E5__MATRIX_ID_SZ 32

`define URAM288E5__NUM_UNIQUE_SELF_ADDR_A    32'h00000418
`define URAM288E5__NUM_UNIQUE_SELF_ADDR_A_SZ 32

`define URAM288E5__NUM_UNIQUE_SELF_ADDR_B    32'h00000419
`define URAM288E5__NUM_UNIQUE_SELF_ADDR_B_SZ 32

`define URAM288E5__NUM_URAM_IN_MATRIX    32'h0000041a
`define URAM288E5__NUM_URAM_IN_MATRIX_SZ 32

`define URAM288E5__OREG_A    32'h0000041b
`define URAM288E5__OREG_A_SZ 40

`define URAM288E5__OREG_B    32'h0000041c
`define URAM288E5__OREG_B_SZ 40

`define URAM288E5__OREG_ECC_A    32'h0000041d
`define URAM288E5__OREG_ECC_A_SZ 40

`define URAM288E5__OREG_ECC_B    32'h0000041e
`define URAM288E5__OREG_ECC_B_SZ 40

`define URAM288E5__PR_SAVE_DATA    32'h0000041f
`define URAM288E5__PR_SAVE_DATA_SZ 40

`define URAM288E5__READ_WIDTH_A    32'h00000420
`define URAM288E5__READ_WIDTH_A_SZ 32

`define URAM288E5__READ_WIDTH_B    32'h00000421
`define URAM288E5__READ_WIDTH_B_SZ 32

`define URAM288E5__REG_CAS_A    32'h00000422
`define URAM288E5__REG_CAS_A_SZ 40

`define URAM288E5__REG_CAS_B    32'h00000423
`define URAM288E5__REG_CAS_B_SZ 40

`define URAM288E5__RST_MODE_A    32'h00000424
`define URAM288E5__RST_MODE_A_SZ 40

`define URAM288E5__RST_MODE_B    32'h00000425
`define URAM288E5__RST_MODE_B_SZ 40

`define URAM288E5__SELF_ADDR_A    32'h00000426
`define URAM288E5__SELF_ADDR_A_SZ 11

`define URAM288E5__SELF_ADDR_B    32'h00000427
`define URAM288E5__SELF_ADDR_B_SZ 11

`define URAM288E5__SELF_MASK_A    32'h00000428
`define URAM288E5__SELF_MASK_A_SZ 11

`define URAM288E5__SELF_MASK_B    32'h00000429
`define URAM288E5__SELF_MASK_B_SZ 11

`define URAM288E5__USE_EXT_CE_A    32'h0000042a
`define URAM288E5__USE_EXT_CE_A_SZ 40

`define URAM288E5__USE_EXT_CE_B    32'h0000042b
`define URAM288E5__USE_EXT_CE_B_SZ 40

`define URAM288E5__WRITE_WIDTH_A    32'h0000042c
`define URAM288E5__WRITE_WIDTH_A_SZ 32

`define URAM288E5__WRITE_WIDTH_B    32'h0000042d
`define URAM288E5__WRITE_WIDTH_B_SZ 32

`endif  // B_URAM288E5_DEFINES_VH