`include "B_X5PLL_INTF_defines.vh"

reg [`X5PLL_INTF_DATA_SZ-1:0] ATTR [0:`X5PLL_INTF_ADDR_N-1];
reg [`X5PLL_INTF__APBCLK_FREQ_SZ-1:0] APBCLK_FREQ_REG = APBCLK_FREQ;
reg [`X5PLL_INTF__DESKEW_SEL_SZ:1] DESKEW_SEL_REG = DESKEW_SEL;
reg [`X5PLL_INTF__DMC_APB_SEL_XPLL_SZ:1] DMC_APB_SEL_XPLL_REG = DMC_APB_SEL_XPLL;
reg [`X5PLL_INTF__DMC_PD_SEL_SZ:1] DMC_PD_SEL_REG = DMC_PD_SEL;
reg [`X5PLL_INTF__RIUCLK_DBLR_BYPASS_SZ:1] RIUCLK_DBLR_BYPASS_REG = RIUCLK_DBLR_BYPASS;
reg [`X5PLL_INTF__RIU_CLK_DBL_DCC_XPLL_SZ-1:0] RIU_CLK_DBL_DCC_XPLL_REG = RIU_CLK_DBL_DCC_XPLL;

initial begin
  ATTR[`X5PLL_INTF__APBCLK_FREQ] = APBCLK_FREQ;
  ATTR[`X5PLL_INTF__DESKEW_SEL] = DESKEW_SEL;
  ATTR[`X5PLL_INTF__DMC_APB_SEL_XPLL] = DMC_APB_SEL_XPLL;
  ATTR[`X5PLL_INTF__DMC_PD_SEL] = DMC_PD_SEL;
  ATTR[`X5PLL_INTF__RIUCLK_DBLR_BYPASS] = RIUCLK_DBLR_BYPASS;
  ATTR[`X5PLL_INTF__RIU_CLK_DBL_DCC_XPLL] = RIU_CLK_DBL_DCC_XPLL;
end

always @(trig_attr) begin
  APBCLK_FREQ_REG = ATTR[`X5PLL_INTF__APBCLK_FREQ];
  DESKEW_SEL_REG = ATTR[`X5PLL_INTF__DESKEW_SEL];
  DMC_APB_SEL_XPLL_REG = ATTR[`X5PLL_INTF__DMC_APB_SEL_XPLL];
  DMC_PD_SEL_REG = ATTR[`X5PLL_INTF__DMC_PD_SEL];
  RIUCLK_DBLR_BYPASS_REG = ATTR[`X5PLL_INTF__RIUCLK_DBLR_BYPASS];
  RIU_CLK_DBL_DCC_XPLL_REG = ATTR[`X5PLL_INTF__RIU_CLK_DBL_DCC_XPLL];
end

// procedures to override, read attribute values

task write_attr;
  input  [`X5PLL_INTF_ADDR_SZ-1:0] addr;
  input  [`X5PLL_INTF_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`X5PLL_INTF_DATA_SZ-1:0] read_attr;
  input  [`X5PLL_INTF_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
