-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : J.PIQUEMAL
--             Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 03/09/2024
--
-- Description : This module top regroup all layer of the SpaceFibrelight IP.
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_lib;
 use phy_plus_lane_lib.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

library interlayer_lib;
use interlayer_lib.all;

entity spacefibre_light_top is
   generic(
      G_VC_NUM                         : integer := 8                              --! Number of virtual channel
      );
   port (
      RST_N                            : in  std_logic;                            --! global reset
      CLK                              : in  std_logic;                            --! Main clock
      CLK_TX                           : out  std_logic;                           --! Clock generated by manufacturer IP
      RST_TXCLK_N                      : out  std_logic;                           --! Reset clock generated by manufacturer IP
      -- CLK HSSL signals
      CLK_REF_N                        : in std_logic;                             --! HSSL dedicated clock
      CLK_REF_P                        : in std_logic;                             --! HSSL dedicated clock
      -- FROM/TO Outside
      TX_POS                           : out std_logic;                            --! Positive LVDS serial data send
      TX_NEG                           : out std_logic;                            --! Negative LVDS serial data send
      RX_POS                           : in  std_logic;                            --! Positive LVDS serial data received
      RX_NEG                           : in  std_logic;                            --! Negative LVDS serial data received
      ----------------------- Data-Link layer signals -----------------------
      -- Discret signals
      AXIS_ARSTN_TX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Active-low asynchronous reset signals for each virtual channel (VC) in the TX path
      AXIS_ACLK_TX_DL                  : in  std_logic_vector(G_VC_NUM downto 0);  --! Clock signals for each VC in the TX path
      AXIS_TREADY_TX_DL                : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates that the data link layer is ready to accept data on each VC
      AXIS_TDATA_TX_DL                 : in  vc_data_array(G_VC_NUM downto 0);     --! Data signals from the network layer to the data link layer for each VC
      AXIS_TUSER_TX_DL                 : in  vc_k_array(G_VC_NUM downto 0);        --! Sideband information (e.g., control or metadata) from the network layer to the data link layer for each VC
      AXIS_TLAST_TX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates the last transfer in a packet/transaction on each VC
      AXIS_TVALID_TX_DL                : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates that valid data is available on the TX data bus for each VC
      AXIS_ARSTN_RX_DL                 : in  std_logic_vector(G_VC_NUM downto 0);  --! Active-low asynchronous reset signals for each VC in the RX path
      AXIS_ACLK_RX_DL                  : in  std_logic_vector(G_VC_NUM downto 0);  --! Clock signals for each VC in the RX path
      AXIS_TREADY_RX_DL                : in  std_logic_vector(G_VC_NUM downto 0);  --! Indicates that the network layer is ready to receive data on each VC
      AXIS_TDATA_RX_DL                 : out vc_data_array(G_VC_NUM downto 0);     --! Data signals from the data link layer to the network layer for each VC
      AXIS_TUSER_RX_DL                 : out vc_k_array(G_VC_NUM downto 0);        --! Sideband information from the data link layer to the network layer for each VC
      AXIS_TLAST_RX_DL                 : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates the last transfer in a packet/transaction on each VC
      AXIS_TVALID_RX_DL                : out std_logic_vector(G_VC_NUM downto 0);  --! Indicates that valid data is available on the RX data bus for each VC
      CURRENT_TIME_SLOT_NW             : in  std_logic_vector(7 downto 0);         --! Current time slot
      -- Paramters signals
      INTERFACE_RESET                  : in  std_logic;                            --! Reset the link and all configuration register of the Data Link layer
      LINK_RESET                       : in  std_logic;                            --! Reset the link
      NACK_RST_EN                      : in  std_logic;                            --! Enable automatic link reset on NACK reception
      NACK_RST_MODE                    : in  std_logic;                            --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
      PAUSE_VC                         : in  std_logic_vector(8 downto 0);         --! Pause the corresponding virtual channel after the end of current transmission
      CONTINUOUS_VC                    : in  std_logic_vector(7 downto 0);         --! Enable the corresponding virtual channel continuous mode
      -- Status signals
      SEQ_NUMBER_TX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in transmission
      SEQ_NUMBER_RX                    : out std_logic_vector(7 downto 0);          --! SEQ_NUMBER in reception
      CREDIT_VC                        : out std_logic_vector(7 downto 0);          --! Indicates if each corresponding far-end input buffer has credit
      INPUT_BUF_OVF_VC                 : out std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates input buffer overflow
      FCT_CREDIT_OVERFLOW              : out std_logic_vector(7 downto 0);          --! Indicates overflow of each corresponding input buffer
      CRC_LONG_ERROR                   : out std_logic;                             --! CRC long error
      CRC_SHORT_ERROR                  : out std_logic;                             --! CRC short error
      FRAME_ERROR                      : out std_logic;                             --! Frame error
      SEQUENCE_ERROR                   : out std_logic;                             --! Sequence error
      FAR_END_LINK_RESET               : out std_logic;                             --! Far-end link reset status
      FRAME_FINISHED                   : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel finished emitting a frame
      FRAME_TX                         : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel is emitting a frame
      DATA_COUNTER_TX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data transmitted in last frame emitted
      DATA_COUNTER_RX                  : out std_logic_vector(6 downto 0);          --! Indicate the number of data received in last frame received
      ACK_COUNTER_TX                   : out std_logic_vector(2 downto 0);          --! ACK counter TX
      NACK_COUNTER_TX                  : out std_logic_vector(2 downto 0);          --! NACK counter TX
      FCT_COUNTER_TX                   : out std_logic_vector(3 downto 0);          --! FCT counter TX
      ACK_COUNTER_RX                   : out std_logic_vector(2 downto 0);          --! ACK counter RX
      NACK_COUNTER_RX                  : out std_logic_vector(2 downto 0);          --! NACK counter RX
      FCT_COUNTER_RX                   : out std_logic_vector(3 downto 0);          --! FCT counter RX
      FULL_COUNTER_RX                  : out std_logic_vector(1 downto 0);          --! FULL counter RX
      RETRY_COUNTER_RX                 : out std_logic_vector(1 downto 0);          --! RETRY counter RX
      CURRENT_TIME_SLOT                : out std_logic_vector(7 downto 0);          --! Current time slot
      RESET_PARAM                      : out std_logic;                             --! Reset parameters register command
      LINK_RST_ASSERTED                : out std_logic;                             --! Link reset status
      NACK_SEQ_NUM                     : out std_logic_vector(7 downto 0);          --! NACK Seq_num received
      ACK_SEQ_NUM                      : out std_logic_vector(7 downto 0);          --! ACK Seq_num received
      DATA_PULSE_RX                    : out std_logic;                             --! Data received pulse signal
      ACK_PULSE_RX                     : out std_logic;                             --! ACK received pulse signal
      NACK_PULSE_RX                    : out std_logic;                             --! NACK received pulse signal
      FCT_PULSE_RX                     : out std_logic;                             --! FCT received pulse signal
      FULL_PULSE_RX                    : out std_logic;                             --! FULL received pulse signal
      RETRY_PULSE_RX                   : out std_logic;                             --! RETRY received pulse signal
      ----------------------- Phy + Lane layer signals -----------------------
      -- -- Interface injector
      ENABLE_INJ                       : in std_logic;                              --! Enable injector command
      DATA_TX_INJ                      : in  std_logic_vector(31 downto 00);        --! Data parallel to be send from injector
      CAPABILITY_TX_INJ                : in  std_logic_vector(07 downto 00);        --! Capability send on TX link in INIT3 control word from injector
      NEW_DATA_TX_INJ                  : in  std_logic;                             --! Flag to write data in FIFO TX from injetor
      VALID_K_CHARAC_TX_INJ            : in  std_logic_vector(03 downto 00);        --! K charachter valid in the 32-bit DATA_TX_INJ vector
      FIFO_TX_FULL_INJ                 : out   std_logic;                           --! Flag full of the FIFO TX to the injector
      LANE_RESET_INJ                   : in  std_logic;                             --! Lane Reset command from Injector
      -- -- Interface spy
      ENABLE_SPY                       : in std_logic;                              --! Enable Spy read command
      FIFO_RX_RD_EN_SPY                : in  std_logic;                             --! FiFo RX read enable flag from the spy
      DATA_RX_SPY                      : out std_logic_vector(31 downto 00);        --! 32-bit Data parallel to be received to the spy
      FIFO_RX_EMPTY_SPY                : out std_logic;                             --! FiFo RX empty flag to the spy
      FIFO_RX_DATA_VALID_SPY           : out std_logic;                             --! FiFo RX data valid flag to the spy
      VALID_K_CHARAC_RX_SPY            : out std_logic_vector(03 downto 00);        --! 4-bit valid K character flags to the spy
      -- Paramter and Status signals
      LANE_START                       : in  std_logic;                             --! Asserts or de-asserts LaneStart for the lane
      AUTOSTART                        : in  std_logic;                             --! Asserts or de-asserts AutoStart for the lane
      LANE_RESET                       : in  std_logic;                             --! Asserts or de-asserts LaneReset for the lane
      PARALLEL_LOOPBACK_EN             : in  std_logic;                             --! Enables or disables the parallel loopback for the lane
      STANDBY_REASON                   : in  std_logic_vector(07 downto 00);        --! In case of error, pauses communication
      NEAR_END_SERIAL_LB_EN            : in  std_logic;                             --! Enables or disables the near-end serial loopback for the lane
      FAR_END_SERIAL_LB_EN             : in  std_logic;                             --! Enables or disables the far-end serial loopback for the lane
      LANE_STATE                       : out std_logic_vector(03 downto 00);        --! Indicates the current state of the Lane Initialization state machine in a lane
      RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);        --! Counter of error detected on the RX link
      RX_ERROR_OVF                     : out std_logic;                             --! Overflow flag of the RX_ERROR_CNT
      LOSS_SIGNAL                      : out std_logic;                             --! Set when no signal is received on RX link
      FAR_END_CAPA                     : out std_logic_vector(07 downto 00);        --! RX Capabilities field (INT3 flags)
      RX_POLARITY                      : out std_logic                              --! Set when the receiver polarity is inverted
   );
end spacefibre_light_top;

architecture rtl of spacefibre_light_top is

   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Modules Declaration -----------------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
   component reset_gen is
      port(
         RST_N                : in  std_logic;     --! global reset
         CLK                  : in  std_logic;     --! General clock
         RST_TX_DONE          : in  std_logic;     --! PLL lock flag
         LANE_RESET           : in  std_logic;     --! LANE RESET command
         INTERNAL_SYNC_RST_N  : out std_logic      --! Internal reset resynchronized on 50MHz internal clock
      );
   end component;

   component data_link is
      generic(
         G_VC_NUM           : integer := 8                                         --! Number of virtual channel
         );
         port(
            RST_N                  : in  std_logic;                                --! global reset
            CLK                    : in  std_logic;                                --! Clock generated by GTY IP
            -- Network layer AXI-Stream TX interface
            AXIS_ARSTN_TX_NW       : in  std_logic_vector(G_VC_NUM downto 0);      --! Active-low asynchronous reset signals for each virtual channel (VC) in the TX path
            AXIS_ACLK_TX_NW        : in  std_logic_vector(G_VC_NUM downto 0);      --! Clock signals for each VC in the TX path
            AXIS_TREADY_TX_DL      : out std_logic_vector(G_VC_NUM downto 0);      --! Indicates that the data link layer is ready to accept data on each VC
            AXIS_TDATA_TX_NW       : in  vc_data_array(G_VC_NUM downto 0);         --! Data signals from the network layer to the data link layer for each VC
            AXIS_TUSER_TX_NW       : in  vc_k_array(G_VC_NUM downto 0);            --! Sideband information (e.g., control or metadata) from the network layer to the data link layer for each VC
            AXIS_TLAST_TX_NW       : in  std_logic_vector(G_VC_NUM downto 0);      --! Indicates the last transfer in a packet/transaction on each VC
            AXIS_TVALID_TX_NW      : in  std_logic_vector(G_VC_NUM downto 0);      --! Indicates that valid data is available on the TX data bus for each VC
            -- Network layer RX interface
            AXIS_ARSTN_RX_NW       : in std_logic_vector(G_VC_NUM downto 0);       --! Active-low asynchronous reset signals for each VC in the RX path
            AXIS_ACLK_RX_NW        : in std_logic_vector(G_VC_NUM downto 0);       --! Clock signals for each VC in the RX path
            AXIS_TREADY_RX_NW      : in  std_logic_vector(G_VC_NUM downto 0);      --! Indicates that the network layer is ready to receive data on each VC
            AXIS_TDATA_RX_DL       : out vc_data_array(G_VC_NUM downto 0);         --! Data signals from the data link layer to the network layer for each VC
            AXIS_TUSER_RX_DL       : out vc_k_array(G_VC_NUM downto 0);            --! Sideband information from the data link layer to the network layer for each VC
            AXIS_TLAST_RX_DL       : out std_logic_vector(G_VC_NUM downto 0);      --! Indicates the last transfer in a packet/transaction on each VC
            AXIS_TVALID_RX_DL      : out std_logic_vector(G_VC_NUM downto 0);      --! Indicates that valid data is available on the RX data bus for each VC
            CURRENT_TIME_SLOT_NW   : in  std_logic_vector(7 downto 0);             --! Current time slot
            -- Lane layer TX interface
            DATA_TX_DL             : out  std_logic_vector(31 downto 00);          --! Data parallel to be send from Data-Link Layer
            CAPABILITY_TX_DL       : out  std_logic_vector(07 downto 00);          --! Capability send on TX link in INIT3 control word
            NEW_DATA_TX_DL         : out  std_logic;                               --! Flag to write data in FIFO TX
            VALID_K_CHARAC_TX_DL   : out  std_logic_vector(03 downto 00);          --! K charachter valid in the 32-bit DATA_TX_DL vector
            FIFO_TX_FULL_PPL       : in   std_logic;                               --! Flag full of the FIFO TX
            -- Lane layer RX interface
            FIFO_RX_RD_EN_DL        : out  std_logic;                              --! Flag to read data in FIFO RX
            DATA_RX_PPL             : in   std_logic_vector(31 downto 00);         --! Data parallel to be received to Data-Link Layer
            FIFO_RX_EMPTY_PPL       : in   std_logic;                              --! Flag EMPTY of the FIFO RX
            FIFO_RX_DATA_VALID_PPL  : in   std_logic;                              --! Flag DATA_VALID of the FIFO RX
            VALID_K_CHARAC_RX_PPL   : in   std_logic_vector(03 downto 00);         --! K charachter valid in the 32-bit DATA_TR_PPL vector
            FAR_END_CAPA_PPL        : in   std_logic_vector(07 downto 00);         --! Capability field receive in INIT3 control word
            LANE_ACTIVE_PPL         : in  std_logic;                               --! Lane Active flag for the DATA Link Layer
            LANE_RESET_DL           : out std_logic;                               --! Lane Reset command
            -- MIB  parameters interface
            INTERFACE_RESET_MIB     : in std_logic;                                --! Reset the link and all configuration register
            LINK_RESET_MIB          : in std_logic;                                --! Reset the link
            NACK_RST_EN_MIB         : in std_logic;                                --! Enable automatic link reset on NACK reception
            NACK_RST_MODE_MIB       : in std_logic;                                --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
            PAUSE_VC_MIB            : in std_logic_vector(G_VC_NUM downto 0);      --! Pause the corresponding virtual channel after the end of current transmission
            CONTINUOUS_VC_MIB       : in std_logic_vector(G_VC_NUM-1 downto 0);    --! Enable the corresponding virtual channel continuous mode
            -- MIB  status interface
            SEQ_NUMBER_TX_DL        : out std_logic_vector(8-1 downto 0);          --! SEQ_NUMBER in transmission
            SEQ_NUMBER_RX_DL        : out std_logic_vector(8-1 downto 0);          --! SEQ_NUMBER in reception
            CREDIT_VC_DL            : out std_logic_vector(G_VC_NUM-1 downto 0);   --! Indicates if each corresponding far-end input buffer has credit
            INPUT_BUF_OVF_VC_DL     : out std_logic_vector(G_VC_NUM-1 downto 0);   --! Indicates input buffer overflow
            FCT_CREDIT_OVERFLOW_DL  : out std_logic_vector(G_VC_NUM-1 downto 0);   --! Indicates overflow of each corresponding input buffer
            CRC_LONG_ERROR_DL       : out std_logic;                               --! CRC long error
            CRC_SHORT_ERROR_DL      : out std_logic;                               --! CRC short error
            FRAME_ERROR_DL          : out std_logic;                               --! Frame error
            SEQUENCE_ERROR_DL       : out std_logic;                               --! Sequence error
            FAR_END_LINK_RESET_DL   : out std_logic;                               --! Far-end link reset status
            FRAME_FINISHED_DL       : out std_logic_vector(G_VC_NUM downto 0);     --! Indicates that corresponding channel finished emitting a frame
            FRAME_TX_DL             : out std_logic_vector(G_VC_NUM downto 0);     --! Indicates that corresponding channel is emitting a frame
            DATA_COUNTER_TX_DL      : out std_logic_vector(6 downto 0);            --! Indicate the number of data transmitted in last frame emitted
            DATA_COUNTER_RX_DL      : out std_logic_vector(6 downto 0);            --! Indicate the number of data received in last frame received
            ACK_COUNTER_TX_DL       : out  std_logic_vector(2 downto 0);           --! ACK counter TX
            NACK_COUNTER_TX_DL      : out  std_logic_vector(2 downto 0);           --! NACK counter TX
            FCT_COUNTER_TX_DL       : out  std_logic_vector(3 downto 0);           --! FCT counter TX
            ACK_COUNTER_RX_DL       : out  std_logic_vector(2 downto 0);           --! ACK counter RX
            NACK_COUNTER_RX_DL      : out  std_logic_vector(2 downto 0);           --! NACK counter RX
            FCT_COUNTER_RX_DL       : out  std_logic_vector(3 downto 0);           --! FCT counter RX
            FULL_COUNTER_RX_DL      : out  std_logic_vector(1 downto 0);           --! FULL counter RX
            RETRY_COUNTER_RX_DL     : out  std_logic_vector(1 downto 0);           --! RETRY counter RX
            CURRENT_TIME_SLOT_DL    : out  std_logic_vector(7 downto 0);           --! Current time slot
            RESET_PARAM_DL          : out std_logic;                               --! Reset configuration parameters control
            LINK_RST_ASSERTED_DL    : out std_logic;                               --! Link has been reseted
            NACK_SEQ_NUM_DL         : out std_logic_vector(7 downto 0);            --! NACK Seq_num received
            ACK_SEQ_NUM_DL          : out std_logic_vector(7 downto 0);            --! ACK Seq_num received
            DATA_PULSE_RX_DL        : out std_logic;                               --! Data received pulse signal
            ACK_PULSE_RX_DL         : out std_logic;                               --! ACK received pulse signal
            NACK_PULSE_RX_DL        : out std_logic;                               --! NACK received pulse signal
            FCT_PULSE_RX_DL         : out std_logic;                               --! FCT received pulse signal
            FULL_PULSE_RX_DL        : out std_logic;                               --! FULL received pulse signal
            RETRY_PULSE_RX_DL       : out std_logic                                --! RETRY received pulse signal
          );
    end component;

    component mux_tx is
      port (
        RST_N                  : in  std_logic;                          --! Global reset
        CLK                    : in  std_logic;                          --! Global clock
        -- Ctrl signal
        ENABLE_INJ             : in std_logic;                           --! Enable injector command
        -- Injector interface
        DATA_TX_INJ            : in  std_logic_vector(31 downto 00);     --! Data parallel to be send from injector
        CAPABILITY_TX_INJ      : in  std_logic_vector(07 downto 00);     --! Capability send on TX link in INIT3 control word from injector
        NEW_DATA_TX_INJ        : in  std_logic;                          --! Flag to write data in FIFO TX from injetor
        VALID_K_CHARAC_TX_INJ  : in  std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TX_INJ vector
        FIFO_TX_FULL_INJ       : out std_logic;                          --! Fifo TX full flag to Injector
        LANE_RESET_INJ         : in  std_logic;                          --! Lane Reset command from Injector
	    	-- Data-Link interface
        DATA_TX_DL             : in  std_logic_vector(31 downto 00);     --! Data parallel to be send from Data-Link Layer
        CAPABILITY_TX_DL       : in  std_logic_vector(07 downto 00);     --! Capability send on TX link in INIT3 control word
        NEW_DATA_TX_DL         : in  std_logic;                          --! Flag to write data in FIFO TX
        VALID_K_CHARAC_TX_DL   : in  std_logic_vector(03 downto 00);     --! K charachter valid in the 32-bit DATA_TX_DL vector
        FIFO_TX_FULL_DL        : out std_logic;                          --! Fifo TX full flag to dl
        LANE_RESET_DL          : in  std_logic;                          --! Lane Reset command from dl
        -- Phy Plus Lane interface
        DATA_TX_MUX            : out  std_logic_vector(31 downto 00);    --! Data parallel
        CAPABILITY_TX_MUX      : out  std_logic_vector(07 downto 00);    --! Capability send on TX link in INIT3 control word
        NEW_DATA_TX_MUX        : out  std_logic;                         --! Flag to write data in FIFO TX
        VALID_K_CHARAC_TX_MUX  : out  std_logic_vector(03 downto 00);    --! K charachter valid in the 32-bit DATA_TX_MUX vector
        FIFO_TX_FULL_PPL       : in   std_logic;                         --! Fifo TX full flag from ppl
        LANE_RESET_MUX         : out  std_logic                          --! Lane Reset command to ppl
  );
   end component;

   component demux_rx is
      port (
        RST_N                  : in  std_logic; --! Global reset
        CLK                    : in  std_logic; --! Global Clock
        -- Ctrl signal
        ENABLE_SPY             : in std_logic;  --! Enable Spy read command
        -- Data-Link interface
        FIFO_RX_RD_EN_DL       : in  std_logic; --! Flag to read data in FIFO RX from Data-Link
        -- SPY interface
        FIFO_RX_RD_EN_SPY      : in  std_logic; --! Flag to read data in FIFO RX from Spy
        -- Phy Plus Lane interface
        FIFO_RX_RD_EN_DEMUX    : out std_logic  --! Flag to read data in FIFO RX to PPL
      );
   end component;

   component phy_plus_lane_64b is
      port(
         RST_N                            : in  std_logic;                       -- global reset
         CLK                              : in  std_logic;                       -- Main clock
         -- Reset_gen interface
         LANE_RESET_PPL_OUT               : out std_logic;
         RST_TXCLK_N                      : in  std_logic;                       -- Synchronous reset on clock generated by GTY PLL
         CLK_TX_OUT                       : out std_logic;                       -- Clock generated by manufacturer IP
         RST_TX_DONE                      : out std_logic;                       -- Up when internal rx reset done
         -- CLK GTY signals
         CLK_REF_N                          : in std_logic;
         CLK_REF_P                          : in std_logic;
         -- FROM Data-link layer
         DATA_TX                          : in  std_logic_vector(31 downto 00);  -- 32-bit Data parallel to be send from Data-Link Layer
         LANE_RESET_DL                    : in  std_logic;                       -- Lane reset command from Data-Link Layer
         CAPABILITY_TX                    : in  std_logic_vector(07 downto 00);  -- Capability field send in INIT3 control word
         NEW_DATA_TX                      : in  std_logic;                       -- Flag new data
         VALID_K_CHARAC_TX                : in  std_logic_vector(03 downto 00);  -- 4-bit valid K character flags from Data-link layer
         FIFO_TX_FULL                     : out std_logic;                       -- FiFo TX full flag

         -- TO Data-link layer
         FIFO_RX_RD_EN                    : in  std_logic;                       -- FiFo RX read enable flag
         DATA_RX                          : out std_logic_vector(31 downto 00);  -- 32-bit Data parallel to be received to Data-Link Layer.
         FIFO_RX_EMPTY                    : out std_logic;                       -- FiFo RX empty flag
         FIFO_RX_DATA_VALID               : out std_logic;                       --! FiFo RX data valid flag
         VALID_K_CHARAC_RX                : out std_logic_vector(03 downto 00);  -- 4-bit valid K character flags to Data-link layer
         FAR_END_CAPA_DL                  : out std_logic_vector(07 downto 00);  -- Capability field receive in INIT3 control word
         LANE_ACTIVE_DL                   : out std_logic;                       -- Lane Active flag for the DATA Link Layer
         -- FROM/TO Outside
         TX_POS                           : out std_logic;                       -- Positive LVDS serial data send
         TX_NEG                           : out std_logic;                       -- Negative LVDS serial data send
         RX_POS                           : in  std_logic;                       -- Positive LVDS serial data received
         RX_NEG                           : in  std_logic;                       -- Negative LVDS serial data received

         -- PARAMETERS and STATUS
         LANE_START                       : in  std_logic;                       -- Asserts or de-asserts LaneStart for the lane
         AUTOSTART                        : in  std_logic;                       -- Asserts or de-asserts AutoStart for the lane
         LANE_RESET                       : in  std_logic;                       -- Asserts or de-asserts LaneReset for the lane
         PARALLEL_LOOPBACK_EN             : in  std_logic;                       -- Enables or disables the parallel loopback for the lane
         STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  -- In case of error, pauses communication
         NEAR_END_SERIAL_LB_EN            : in  std_logic;                       -- Enables or disables the near-end serial loopback for the lane
         FAR_END_SERIAL_LB_EN             : in  std_logic;                       -- Enables or disables the far-end serial loopback for the lane

         LANE_STATE                       : out std_logic_vector(03 downto 00);  -- Indicates the current state of the Lane Initialization state machine in a lane
         RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  -- Counter of error detected on the RX link
         RX_ERROR_OVF                     : out std_logic;                       -- Overflow flag of the RX_ERROR_CNT
         LOSS_SIGNAL                      : out std_logic;                       -- Set when no signal is received on RX link
         FAR_END_CAPA                     : out std_logic_vector(07 downto 00);  -- Capabilities field (INT3 flags)
         RX_POLARITY                      : out std_logic                        -- Set when the receiver polarity is inverted
      );
   end component;
   component mib_data_link is
      generic(
          G_VC_NUM               : integer := 8                                --! Number of virtual channel
         );
        port (
          -- MIB parameters interface TOP
          INTERFACE_RESET         : in  std_logic;                             --! Reset the link and all configuration register of the Data Link layer from the TOP
          LINK_RESET              : in  std_logic;                             --! Reset the link from the TOP
          NACK_RST_EN             : in  std_logic;                             --! Enable automatic link reset on NACK reception from the TOP
          NACK_RST_MODE           : in  std_logic;                             --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception from the TOP
          PAUSE_VC                : in  std_logic_vector(G_VC_NUM downto 0);   --! Pause the corresponding virtual channel after the end of current transmission from the TOP
          CONTINUOUS_VC           : in  std_logic_vector(G_VC_NUM-1 downto 0); --! Enable the corresponding virtual channel continuous mode from the TOP
          -- MIB parameters interface Data-link
          INTERFACE_RESET_DL      : out std_logic;                             --! Reset the link and all configuration register of the Data Link layer to DL
          LINK_RESET_DL           : out std_logic;                             --! Reset the link to DL
          NACK_RST_EN_DL          : out std_logic;                             --! Enable automatic link reset on NACK reception to DL
          NACK_RST_MODE_DL        : out std_logic;                             --! Up for instant link reset on NACK reception, down for link reset at the end of current received frame on NACK reception to DL
          PAUSE_VC_DL             : out std_logic_vector(G_VC_NUM downto 0);   --! Pause the corresponding virtual channel after the end of current transmission to DL
          CONTINUOUS_VC_DL        : out std_logic_vector(G_VC_NUM-1 downto 0); --! Enable the corresponding virtual channel continuous mode to DL
          -- MIB status interface Data-link
          SEQ_NUMBER_TX_DL        : in  std_logic_vector(G_VC_NUM-1 downto 0); --! SEQ_NUMBER in transmission from DL
          SEQ_NUMBER_RX_DL        : in  std_logic_vector(G_VC_NUM-1 downto 0); --! SEQ_NUMBER in reception from DL
          CREDIT_VC_DL            : in  std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates if each corresponding far-end input buffer has credit from DL
          INPUT_BUF_OVF_VC_DL     : in  std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates input buffer overflow from DL
          FCT_CREDIT_OVERFLOW_DL  : in  std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates overflow of each corresponding input buffer from DL
          CRC_LONG_ERROR_DL       : in  std_logic;                             --! CRC long error from DL
          CRC_SHORT_ERROR_DL      : in  std_logic;                             --! CRC short error from DL
          FRAME_ERROR_DL          : in  std_logic;                             --! Frame error from DL
          SEQUENCE_ERROR_DL       : in  std_logic;                             --! Sequence error from DL
          FAR_END_LINK_RESET_DL   : in  std_logic;                             --! Far-end link reset status from DL
          FRAME_FINISHED_DL       : in  std_logic_vector(G_VC_NUM downto 0);   --! Indicates that corresponding channel finished emitting a frame from DL
          FRAME_TX_DL             : in  std_logic_vector(G_VC_NUM downto 0);   --! Indicates that corresponding channel is emitting a frame from DL
          DATA_COUNTER_TX_DL      : in  std_logic_vector(6 downto 0);          --! Indicate the number of data transmitted in last frame emitted from DL
          DATA_COUNTER_RX_DL      : in  std_logic_vector(6 downto 0);          --! Indicate the number of data received in last frame received from DL
          ACK_COUNTER_TX_DL       : in  std_logic_vector(2 downto 0);          --! ACK counter TX from DL
          NACK_COUNTER_TX_DL      : in  std_logic_vector(2 downto 0);          --! NACK counter TX from DL
          FCT_COUNTER_TX_DL       : in  std_logic_vector(3 downto 0);          --! FCT counter TX from DL
          ACK_COUNTER_RX_DL       : in  std_logic_vector(2 downto 0);          --! ACK counter RX from DL
          NACK_COUNTER_RX_DL      : in  std_logic_vector(2 downto 0);          --! NACK counter RX from DL
          FCT_COUNTER_RX_DL       : in  std_logic_vector(3 downto 0);          --! FCT counter RX from DL
          FULL_COUNTER_RX_DL      : in  std_logic_vector(1 downto 0);          --! FULL counter RX from DL
          RETRY_COUNTER_RX_DL     : in  std_logic_vector(1 downto 0);          --! RETRY counter RX from DL
          CURRENT_TIME_SLOT_DL    : in  std_logic_vector(G_VC_NUM-1 downto 0); --! Current time slot from DL
          RESET_PARAM_DL          : in  std_logic;                             --! Reset configuration parameters control from DL
          LINK_RST_ASSERTED_DL    : in  std_logic;                             --! Link has been reseted from DL
          NACK_SEQ_NUM_DL         : in std_logic_vector(7 downto 0);           --! NACK Seq_num received from DL
          ACK_SEQ_NUM_DL          : in std_logic_vector(7 downto 0);           --! ACK Seq_num received from DL
          DATA_PULSE_RX_DL        : in std_logic;                              --! Data received pulse signal from DL
          ACK_PULSE_RX_DL         : in std_logic;                              --! ACK received pulse signal from DL
          NACK_PULSE_RX_DL        : in std_logic;                              --! NACK received pulse signal from DL
          FCT_PULSE_RX_DL         : in std_logic;                              --! FCT received pulse signal from DL
          FULL_PULSE_RX_DL        : in std_logic;                              --! FULL received pulse signal from DL
          RETRY_PULSE_RX_DL       : in std_logic;                              --! RETRY received pulse signal from DL
          -- MIB status interface TOP
          SEQ_NUMBER_TX           : out std_logic_vector(G_VC_NUM-1 downto 0); --! SEQ_NUMBER in transmission to the TOP
          SEQ_NUMBER_RX           : out std_logic_vector(G_VC_NUM-1 downto 0); --! SEQ_NUMBER in reception to the TOP
          CREDIT_VC               : out std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates if each corresponding far-end input buffer has credit to the TOP
          INPUT_BUF_OVF_VC        : out std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates input buffer overflow to the TOP
          FCT_CREDIT_OVERFLOW     : out std_logic_vector(G_VC_NUM-1 downto 0); --! Indicates overflow of each corresponding input buffer to the TOP
          CRC_LONG_ERROR          : out std_logic;                             --! CRC long error to the TOP
          CRC_SHORT_ERROR         : out std_logic;                             --! CRC short error to the TOP
          FRAME_ERROR             : out std_logic;                             --! Frame error to the TOP
          SEQUENCE_ERROR          : out std_logic;                             --! Sequence error to the TOP
          FAR_END_LINK_RESET      : out std_logic;                             --! Far-end link reset status to the TOP
          FRAME_FINISHED          : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel finished emitting a frame to the TOP
          FRAME_TX                : out std_logic_vector(8 downto 0);          --! Indicates that corresponding channel is emitting a frame to the TOP
          DATA_COUNTER_TX         : out std_logic_vector(6 downto 0);          --! Indicate the number of data transmitted in last frame emitted to the TOP
          DATA_COUNTER_RX         : out std_logic_vector(6 downto 0);          --! Indicate the number of data received in last frame received to the TOP
          ACK_COUNTER_TX          : out std_logic_vector(2 downto 0);          --! ACK counter TX to the TOP
          NACK_COUNTER_TX         : out std_logic_vector(2 downto 0);          --! NACK counter TX to the TOP
          FCT_COUNTER_TX          : out std_logic_vector(3 downto 0);          --! FCT counter TX to the TOP
          ACK_COUNTER_RX          : out std_logic_vector(2 downto 0);          --! ACK counter RX to the TOP
          NACK_COUNTER_RX         : out std_logic_vector(2 downto 0);          --! NACK counter RX to the TOP
          FCT_COUNTER_RX          : out std_logic_vector(3 downto 0);          --! FCT counter RX to the TOP
          FULL_COUNTER_RX         : out std_logic_vector(1 downto 0);          --! FULL counter RX to the TOP
          RETRY_COUNTER_RX        : out std_logic_vector(1 downto 0);          --! RETRY counter RX to the TOP
          CURRENT_TIME_SLOT       : out std_logic_vector(G_VC_NUM-1 downto 0); --! Current time slot to the TOP
          RESET_PARAM             : out std_logic;                             --! Reset configuration parameters control to the TOP
          LINK_RST_ASSERTED       : out std_logic;                             --! Link has been reseted to the TOP
          NACK_SEQ_NUM            : out std_logic_vector(7 downto 0);          --! NACK Seq_num received to the TOP
          ACK_SEQ_NUM             : out std_logic_vector(7 downto 0);          --! ACK Seq_num received to the TOP
          DATA_PULSE_RX           : out std_logic;                             --! Data received pulse signal to the TOP
          ACK_PULSE_RX            : out std_logic;                             --! ACK received pulse signal to the TOP
          NACK_PULSE_RX           : out std_logic;                             --! NACK received pulse signal to the TOP
          FCT_PULSE_RX            : out std_logic;                             --! FCT received pulse signal to the TOP
          FULL_PULSE_RX           : out std_logic;                             --! FULL received pulse signal to the TOP
          RETRY_PULSE_RX          : out std_logic                              --! RETRY received pulse signal to the TOP
   );
   end component;

   component mib_phy_plus_lane is
      port(
         -- Parameters From USERAPP/TOP
         LANE_START                       : in  std_logic;                       -- Asserts or de-asserts LaneStart for the lane
         AUTOSTART                        : in  std_logic;                       -- Asserts or de-asserts AutoStart for the lane
         LANE_RESET                       : in  std_logic;                       -- Asserts or de-asserts LaneReset for the lane
         PARALLEL_LOOPBACK_EN             : in  std_logic;                       -- Enables or disables the parallel loopback for the lane.
         STANDBY_REASON                   : in  std_logic_vector(07 downto 00);  -- In case of error, pauses communication.
         NEAR_END_SERIAL_LB_EN            : in  std_logic;                       -- Enables or disables the near-end serial loopback for the lane
         FAR_END_SERIAL_LB_EN             : in  std_logic;                       -- Enables or disables the far-end serial loopback for the lane
         -- Status To USERAPP/TOP
         LANE_STATE                       : out std_logic_vector(03 downto 00);  -- Indicates the current state of the Lane Initialization state machine in a lane
         RX_ERROR_CNT                     : out std_logic_vector(07 downto 00);  -- Counter of error detected on the RX link
         RX_ERROR_OVF                     : out std_logic;                       -- Overflow flag of the RX_ERROR_CNT
         LOSS_SIGNAL                      : out std_logic;                       -- Set when no signal is received on RX link
         FAR_END_CAPA                     : out std_logic_vector(07 downto 00);  -- Capabilities field (INT3 flags)
         RX_POLARITY                      : out std_logic;                       -- Set when the receiver polarity is inverted
         -- Parameters to Module PHY+LANE
         LANE_START_TO_MOD                : out std_logic;                       -- Asserts or de-asserts LaneStart for the lane
         AUTOSTART_TO_MOD                 : out std_logic;                       -- Asserts or de-asserts AutoStart for the lane
         LANE_RESET_TO_MOD                : out std_logic;                       -- Asserts or de-asserts LaneReset for the lane
         PARALLEL_LOOPBACK_EN_TO_MOD      : out std_logic;                       -- Enables or disables the parallel loopback for the lane
         STANDBY_REASON_TO_MOD            : out std_logic_vector(07 downto 00);  -- In case of error, pauses communication
         NEAR_END_SERIAL_LB_EN_TO_MOD     : out std_logic;                       -- Enables or disables the near-end serial loopback for the lane
         FAR_END_SERIAL_LB_EN_TO_MOD      : out std_logic;                       -- Enables or disables the far-end serial loopback for the lane
         -- Status from Module PHY+LANE
         LANE_STATE_FROM_MOD              : in  std_logic_vector(03 downto 00);  -- Indicates the current state of the Lane Initialization state machine in a lane
         RX_ERROR_CNT_FROM_MOD            : in  std_logic_vector(07 downto 00);  -- Counter of error detected on the RX link
         RX_ERROR_OVF_FROM_MOD            : in  std_logic;                       -- Overflow flag of the RX_ERROR_CNT
         LOSS_SIGNAL_FROM_MOD             : in  std_logic;                       -- Set when no signal is received on RX link
         FAR_END_CAPA_FROM_MOD            : in  std_logic_vector(07 downto 00);  -- Capabilities field (INT3 flags)
         RX_POLARITY_FROM_MOD             : in  std_logic                        -- Set when the receiver polarity is inverted
      );
   end component;

   ----------------------------------------------------------------------------------------------------------------------------------------
   -------------------------------------------------------- Internal signals declaration --------------------------------------------------
   ----------------------------------------------------------------------------------------------------------------------------------------
   -- Reset generator internal signals
   signal rst_sync_gty_n                     : std_logic;                        --! Synchronous reset on clock generated by GTY PLL
   -- phy_plus_lane internal signals
   signal clk_tx_i                           : std_logic;                        --! Clock generated by PLL of the manufacturer IP
   signal rst_tx_done                        : std_logic;                         --! Up when internal rx reset done
   signal lane_reset_ppl_out                 : std_logic;
   -- DATA-LINK // Phy plus Lane interface TX signals
   signal data_tx_dl             : std_logic_vector(31 downto 0);  -- Data parallel to be send from Data-Link Layer
   signal capability_tx_dl       : std_logic_vector(7 downto 0);   -- Capability send on TX link in INIT3 control word
   signal new_data_tx_dl         : std_logic;                      -- Flag to write data in FIFO TX
   signal valid_k_charac_tx_dl   : std_logic_vector(3 downto 0);   -- K character valid in the 32-bit DATA_TX_DL vector
   signal fifo_tx_full_mux       : std_logic;                      -- Flag full of the FIFO TX
   -- DATA-LINK // Phy plus Lane interface TX signals
   signal fifo_rx_rd_en_dl       : std_logic;                      -- Flag to read data in FIFO RX
   signal data_rx_ppl            : std_logic_vector(31 downto 0);  -- Data parallel to be received to Data-Link Layer
   signal fifo_rx_empty_ppl      : std_logic;                      -- Flag EMPTY of the FIFO RX
   signal fifo_rx_data_valid_ppl : std_logic;                      -- Flag DATA_VALID of the FIFO RX
   signal valid_k_charac_rx_ppl  : std_logic_vector(3 downto 0);   -- K character valid in the 32-bit DATA_TR_PPL vector
   signal far_end_capa_ppl       : std_logic_vector(7 downto 0);   -- Capability field receive in INIT3 control word
   signal far_end_capa_dl_ppl    : std_logic_vector(7 downto 0);   -- Capability field receive in INIT3 control word
   signal lane_active_ppl        : std_logic;                      -- Lane Active flag for the DATA Link Layer
   signal lane_reset_dl          : std_logic;                      -- Lane Reset flag for the Data Link Layer
   -- MIB phy_plus_lane internal signals
   signal lane_start_ppl                     : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal autostart_ppl                      : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal lane_reset_ppl                     : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal parallel_loopback_en_ppl           : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal standby_reason_ppl                 : std_logic_vector(07 downto 00);   --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal near_end_serial_lb_en_ppl          : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal far_end_serial_lb_en_ppl           : std_logic;                        --! Parameter signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal lane_state_ppl                     : std_logic_vector(03 downto 00);   --! Status signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal rx_error_cnt_ppl                   : std_logic_vector(07 downto 00);   --! Status signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal rx_error_ovf_ppl                   : std_logic;                        --! Status signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal loss_signal_ppl                    : std_logic;                        --! Status signal between MIB_phy_plus_lane and phy_plus_lane modules
   signal rx_polarity_ppl                    : std_logic;                        --! Status signal between MIB_phy_plus_lane and phy_plus_lane modules
   -- MIB data_link internal signals
   signal interface_reset_dl                 : std_logic;
   signal link_reset_dl                      : std_logic;
   signal nack_rst_en_dl                     : std_logic;
   signal nack_rst_mode_dl                   : std_logic;
   signal pause_vc_dl                        : std_logic_vector(G_VC_NUM downto 0);
   signal continuous_vc_dl                   : std_logic_vector(G_VC_NUM-1 downto 0);
   signal seq_number_tx_dl                   : std_logic_vector(G_VC_NUM-1 downto 0);
   signal seq_number_rx_dl                   : std_logic_vector(G_VC_NUM-1 downto 0);
   signal credit_vc_dl                       : std_logic_vector(G_VC_NUM-1 downto 0);
   signal input_buf_ovf_vc_dl                : std_logic_vector(G_VC_NUM-1 downto 0);
   signal fct_credit_overflow_dl             : std_logic_vector(G_VC_NUM-1 downto 0);
   signal crc_long_error_dl                  : std_logic;
   signal crc_short_error_dl                 : std_logic;
   signal frame_error_dl                     : std_logic;
   signal sequence_error_dl                  : std_logic;
   signal far_end_link_reset_dl              : std_logic;
   signal frame_finished_dl                  : std_logic_vector(G_VC_NUM downto 0);
   signal frame_tx_dl                        : std_logic_vector(G_VC_NUM downto 0);
   signal data_counter_tx_dl                 : std_logic_vector(6 downto 0);
   signal data_counter_rx_dl                 : std_logic_vector(6 downto 0);
   signal ack_counter_tx_dl                  : std_logic_vector(2 downto 0);
   signal nack_counter_tx_dl                 : std_logic_vector(2 downto 0);
   signal fct_counter_tx_dl                  : std_logic_vector(3 downto 0);
   signal ack_counter_rx_dl                  : std_logic_vector(2 downto 0);
   signal nack_counter_rx_dl                 : std_logic_vector(2 downto 0);
   signal fct_counter_rx_dl                  : std_logic_vector(3 downto 0);
   signal full_counter_rx_dl                 : std_logic_vector(1 downto 0);
   signal retry_counter_rx_dl                : std_logic_vector(1 downto 0);
   signal current_time_slot_dl               : std_logic_vector(G_VC_NUM-1 downto 0);
   signal reset_param_dl                     : std_logic;
   signal link_rst_asserted_dl               : std_logic;
   signal nack_seq_num_dl                    : std_logic_vector(7 downto 0);
   signal ack_seq_num_dl                     : std_logic_vector(7 downto 0);
   signal data_pulse_rx_dl                   : std_logic;
   signal ack_pulse_rx_dl                    : std_logic;
   signal nack_pulse_rx_dl                   : std_logic;
   signal fct_pulse_rx_dl                    : std_logic;
   signal full_pulse_rx_dl                   : std_logic;
   signal retry_pulse_rx_dl                  : std_logic;
   -- Mux // Phy plus Lane interface TX signals
   signal data_tx_mux                        : std_logic_vector(31 downto 00);
   signal capability_tx_mux                  : std_logic_vector(07 downto 00);
   signal new_data_tx_mux                    : std_logic;
   signal valid_k_charac_tx_mux              : std_logic_vector(03 downto 00);
   signal fifo_tx_full_ppl                   : std_logic;
   signal lane_reset_mux                     : std_logic;
   -- Demux // Phy plus Lane interface TX signals
   signal fifo_rx_rd_en_demux                : std_logic;

begin
   ------------------------------------------------------------------------------------------------------------------
   -------------------------------------------- Reset generator modules ---------------------------------------------
   ------------------------------------------------------------------------------------------------------------------
   inst_reset_sync_clk_from_GTY : reset_gen
   port map(
      RST_N               => RST_N,
      CLK                 => clk_tx_i,
      RST_TX_DONE         => rst_tx_done,
      LANE_RESET          => lane_reset_ppl_out,
      INTERNAL_SYNC_RST_N => rst_sync_gty_n
   );
   -----------------------------------------------------------------------------------------------------------------
   ---------------------------------------------- DATA-LINK layer modules ---------------------------------------------
   ------------------------------------------------------------------------------------------------------------------
   inst_data_link : data_link
   generic map (
      G_VC_NUM => G_VC_NUM
   )
   Port map (
      CLK                      => CLK,
      RST_N                    => RST_N,
       -- Network layer AXI-Stream TX interface
       AXIS_ARSTN_TX_NW        => AXIS_ARSTN_TX_DL,
       AXIS_ACLK_TX_NW         => AXIS_ACLK_TX_DL,
       AXIS_TREADY_TX_DL       => AXIS_TREADY_TX_DL,
       AXIS_TDATA_TX_NW        => AXIS_TDATA_TX_DL,
       AXIS_TUSER_TX_NW        => AXIS_TUSER_TX_DL,
       AXIS_TLAST_TX_NW        => AXIS_TLAST_TX_DL,
       AXIS_TVALID_TX_NW       => AXIS_TVALID_TX_DL,
       -- Network layer RX interface
       AXIS_ARSTN_RX_NW        => AXIS_ARSTN_RX_DL,
       AXIS_ACLK_RX_NW         => AXIS_ACLK_RX_DL,
       AXIS_TREADY_RX_NW       => AXIS_TREADY_RX_DL,
       AXIS_TDATA_RX_DL        => AXIS_TDATA_RX_DL,
       AXIS_TUSER_RX_DL        => AXIS_TUSER_RX_DL,
       AXIS_TLAST_RX_DL        => AXIS_TLAST_RX_DL,
       AXIS_TVALID_RX_DL       => AXIS_TVALID_RX_DL,
       CURRENT_TIME_SLOT_NW    => CURRENT_TIME_SLOT_NW,
       -- Lane layer TX interface
       DATA_TX_DL              =>  data_tx_dl,
       CAPABILITY_TX_DL        =>  capability_tx_dl,
       NEW_DATA_TX_DL          =>  new_data_tx_dl,
       VALID_K_CHARAC_TX_DL    =>  valid_k_charac_tx_dl,
       FIFO_TX_FULL_PPL        =>  fifo_tx_full_mux,
       -- Lane layer RX interface
       FIFO_RX_RD_EN_DL        => fifo_rx_rd_en_dl,
       DATA_RX_PPL             => data_rx_ppl,
       FIFO_RX_EMPTY_PPL       => fifo_rx_empty_ppl,
       FIFO_RX_DATA_VALID_PPL  => fifo_rx_data_valid_ppl,
       VALID_K_CHARAC_RX_PPL   => valid_k_charac_rx_ppl,
       FAR_END_CAPA_PPL        => far_end_capa_dl_ppl,
       LANE_ACTIVE_PPL         => lane_active_ppl,
       LANE_RESET_DL           => lane_reset_dl,
       -- MIB parameters interface
       INTERFACE_RESET_MIB     => interface_reset_dl,
       LINK_RESET_MIB          => link_reset_dl,
       NACK_RST_EN_MIB         => nack_rst_en_dl,
       NACK_RST_MODE_MIB       => nack_rst_mode_dl,
       PAUSE_VC_MIB            => pause_vc_dl,
       CONTINUOUS_VC_MIB       => continuous_vc_dl,
       -- MIB status interface
       SEQ_NUMBER_TX_DL        => seq_number_tx_dl,
       SEQ_NUMBER_RX_DL        => seq_number_rx_dl,
       CREDIT_VC_DL            => credit_vc_dl,
       INPUT_BUF_OVF_VC_DL     => input_buf_ovf_vc_dl,
       FCT_CREDIT_OVERFLOW_DL  => fct_credit_overflow_dl,
       CRC_LONG_ERROR_DL       => crc_long_error_dl,
       CRC_SHORT_ERROR_DL      => crc_short_error_dl,
       FRAME_ERROR_DL          => frame_error_dl,
       SEQUENCE_ERROR_DL       => sequence_error_dl,
       FAR_END_LINK_RESET_DL   => far_end_link_reset_dl,
       FRAME_FINISHED_DL       => frame_finished_dl,
       FRAME_TX_DL             => frame_tx_dl,
       DATA_COUNTER_TX_DL      => data_counter_tx_dl,
       DATA_COUNTER_RX_DL      => data_counter_rx_dl,
       ACK_COUNTER_TX_DL       => ack_counter_tx_dl,
       NACK_COUNTER_TX_DL      => nack_counter_tx_dl,
       FCT_COUNTER_TX_DL       => fct_counter_tx_dl,
       ACK_COUNTER_RX_DL       => ack_counter_rx_dl,
       NACK_COUNTER_RX_DL      => nack_counter_rx_dl,
       FCT_COUNTER_RX_DL       => fct_counter_rx_dl,
       FULL_COUNTER_RX_DL      => full_counter_rx_dl,
       RETRY_COUNTER_RX_DL     => retry_counter_rx_dl,
       CURRENT_TIME_SLOT_DL    => current_time_slot_dl,
       RESET_PARAM_DL          => reset_param_dl,
       LINK_RST_ASSERTED_DL    => link_rst_asserted_dl,
       NACK_SEQ_NUM_DL         => nack_seq_num_dl,
       ACK_SEQ_NUM_DL          => ack_seq_num_dl,
       DATA_PULSE_RX_DL        => data_pulse_rx_dl,
       ACK_PULSE_RX_DL         => ack_pulse_rx_dl,
       NACK_PULSE_RX_DL        => nack_pulse_rx_dl,
       FCT_PULSE_RX_DL         => fct_pulse_rx_dl,
       FULL_PULSE_RX_DL        => full_pulse_rx_dl,
       RETRY_PULSE_RX_DL       => retry_pulse_rx_dl
   );

   inst_mib_data_link : mib_data_link
      generic map (
         G_VC_NUM => G_VC_NUM
      )
      Port map (
         -- MIB parameters interface Lane
         INTERFACE_RESET     => INTERFACE_RESET,
         LINK_RESET          => LINK_RESET,
         NACK_RST_EN         => NACK_RST_EN,
         NACK_RST_MODE       => NACK_RST_MODE,
         PAUSE_VC            => PAUSE_VC,
         CONTINUOUS_VC       => CONTINUOUS_VC,
         -- MIB parameters interface Data-link
         INTERFACE_RESET_DL  => interface_reset_dl,
         LINK_RESET_DL       => link_reset_dl,
         NACK_RST_EN_DL      => nack_rst_en_dl,
         NACK_RST_MODE_DL    => nack_rst_mode_dl,
         PAUSE_VC_DL         => pause_vc_dl,
         CONTINUOUS_VC_DL    => continuous_vc_dl,
         -- MIB status interface Data-link
         SEQ_NUMBER_TX_DL    => seq_number_tx_dl,
         SEQ_NUMBER_RX_DL    => seq_number_rx_dl,
         CREDIT_VC_DL        => credit_vc_dl,
         INPUT_BUF_OVF_VC_DL     => input_buf_ovf_vc_dl,
         FCT_CREDIT_OVERFLOW_DL => fct_credit_overflow_dl,
         CRC_LONG_ERROR_DL   => crc_long_error_dl,
         CRC_SHORT_ERROR_DL  => crc_short_error_dl,
         FRAME_ERROR_DL      => frame_error_dl,
         SEQUENCE_ERROR_DL   => sequence_error_dl,
         FAR_END_LINK_RESET_DL => far_end_link_reset_dl,
         FRAME_FINISHED_DL   => frame_finished_dl,
         FRAME_TX_DL         => frame_tx_dl,
         DATA_COUNTER_TX_DL  => data_counter_tx_dl,
         DATA_COUNTER_RX_DL  => data_counter_rx_dl,
         ACK_COUNTER_TX_DL   => ack_counter_tx_dl,
         NACK_COUNTER_TX_DL  => nack_counter_tx_dl,
         FCT_COUNTER_TX_DL   => fct_counter_tx_dl,
         ACK_COUNTER_RX_DL   => ack_counter_rx_dl,
         NACK_COUNTER_RX_DL  => nack_counter_rx_dl,
         FCT_COUNTER_RX_DL   => fct_counter_rx_dl,
         FULL_COUNTER_RX_DL  => full_counter_rx_dl,
         RETRY_COUNTER_RX_DL => retry_counter_rx_dl,
         CURRENT_TIME_SLOT_DL => current_time_slot_dl,
         RESET_PARAM_DL       => reset_param_dl,
         LINK_RST_ASSERTED_DL => link_rst_asserted_dl,
         NACK_SEQ_NUM_DL      => nack_seq_num_dl,
         ACK_SEQ_NUM_DL       => ack_seq_num_dl,
         DATA_PULSE_RX_DL     => data_pulse_rx_dl,
         ACK_PULSE_RX_DL      => ack_pulse_rx_dl,
         NACK_PULSE_RX_DL     => nack_pulse_rx_dl,
         FCT_PULSE_RX_DL      => fct_pulse_rx_dl,
         FULL_PULSE_RX_DL     => full_pulse_rx_dl,
         RETRY_PULSE_RX_DL    => retry_pulse_rx_dl,
         -- MIB status interface Lane
         SEQ_NUMBER_TX       => SEQ_NUMBER_TX,
         SEQ_NUMBER_RX       => SEQ_NUMBER_RX,
         CREDIT_VC           => CREDIT_VC,
         INPUT_BUF_OVF_VC    => INPUT_BUF_OVF_VC,
         FCT_CREDIT_OVERFLOW => FCT_CREDIT_OVERFLOW,
         CRC_LONG_ERROR      => CRC_LONG_ERROR,
         CRC_SHORT_ERROR     => CRC_SHORT_ERROR,
         FRAME_ERROR         => FRAME_ERROR,
         SEQUENCE_ERROR      => SEQUENCE_ERROR,
         FAR_END_LINK_RESET  => FAR_END_LINK_RESET,
         FRAME_FINISHED      => FRAME_FINISHED,
         FRAME_TX            => FRAME_TX,
         DATA_COUNTER_TX     => DATA_COUNTER_TX,
         DATA_COUNTER_RX     => DATA_COUNTER_RX,
         ACK_COUNTER_TX      => ACK_COUNTER_TX,
         NACK_COUNTER_TX     => NACK_COUNTER_TX,
         FCT_COUNTER_TX      => FCT_COUNTER_TX,
         ACK_COUNTER_RX      => ACK_COUNTER_RX,
         NACK_COUNTER_RX     => NACK_COUNTER_RX,
         FCT_COUNTER_RX      => FCT_COUNTER_RX,
         FULL_COUNTER_RX     => FULL_COUNTER_RX,
         RETRY_COUNTER_RX    => RETRY_COUNTER_RX,
         CURRENT_TIME_SLOT   => CURRENT_TIME_SLOT,
         RESET_PARAM         => RESET_PARAM,
         LINK_RST_ASSERTED   => LINK_RST_ASSERTED,
         NACK_SEQ_NUM        => NACK_SEQ_NUM,
         ACK_SEQ_NUM         => ACK_SEQ_NUM,
         DATA_PULSE_RX       => DATA_PULSE_RX,
         ACK_PULSE_RX        => ACK_PULSE_RX,
         NACK_PULSE_RX       => NACK_PULSE_RX,
         FCT_PULSE_RX        => FCT_PULSE_RX,
         FULL_PULSE_RX       => FULL_PULSE_RX,
         RETRY_PULSE_RX      => RETRY_PULSE_RX
      );
   -----------------------------------------------------------------------------------------------------------------
   ----------------------------------------------- Inter Layer modules ---------------------------------------------
   -----------------------------------------------------------------------------------------------------------------
   ---------------------------------------------------------
   -----                     Assignements              -----
   ---------------------------------------------------------
   DATA_RX_SPY            <= data_rx_ppl;
   FIFO_RX_EMPTY_SPY      <= fifo_rx_empty_ppl;
   FIFO_RX_DATA_VALID_SPY <= fifo_rx_data_valid_ppl;
   VALID_K_CHARAC_RX_SPY  <= valid_k_charac_rx_ppl;
   ---------------------------------------------------------
   -----                     Instantiation             -----
   ---------------------------------------------------------
   inst_mux_tx: mux_tx
      port map(
        RST_N                  => RST_N,
        CLK                    => CLK,
        -- Ctrl signal
        ENABLE_INJ             => ENABLE_INJ,
        -- Injector interface
        DATA_TX_INJ            =>  DATA_TX_INJ,
        CAPABILITY_TX_INJ      =>  CAPABILITY_TX_INJ,
        NEW_DATA_TX_INJ        =>  NEW_DATA_TX_INJ,
        VALID_K_CHARAC_TX_INJ  =>  VALID_K_CHARAC_TX_INJ,
        FIFO_TX_FULL_INJ       =>  FIFO_TX_FULL_INJ,
        LANE_RESET_INJ         =>  LANE_RESET_INJ,
          -- Data-Link interfa
        DATA_TX_DL             => data_tx_dl,
        CAPABILITY_TX_DL       => capability_tx_dl,
        NEW_DATA_TX_DL         => new_data_tx_dl,
        VALID_K_CHARAC_TX_DL   => valid_k_charac_tx_dl,
        FIFO_TX_FULL_DL        => fifo_tx_full_mux,
        LANE_RESET_DL          => lane_reset_dl,
        -- Phy Plus Lane interf
        DATA_TX_MUX            => data_tx_mux,
        CAPABILITY_TX_MUX      => capability_tx_mux,
        NEW_DATA_TX_MUX        => new_data_tx_mux,
        VALID_K_CHARAC_TX_MUX  => valid_k_charac_tx_mux,
        FIFO_TX_FULL_PPL       => fifo_tx_full_ppl,
        LANE_RESET_MUX         => lane_reset_mux
      );
   inst_demux_rx: demux_rx
      port map (
        RST_N                  => RST_N,
        CLK                    => CLK,
        -- Ctrl signal
        ENABLE_SPY             => ENABLE_SPY,
        -- Data-Link Interface
        FIFO_RX_RD_EN_DL       => fifo_rx_rd_en_dl,
        -- SPY interface
        FIFO_RX_RD_EN_SPY      => FIFO_RX_RD_EN_SPY,
        -- Phy Plus Lane int
        FIFO_RX_RD_EN_DEMUX    => fifo_rx_rd_en_demux
      );
   -----------------------------------------------------------------------------------------------------------------
   ---------------------------------------------- PHY_PLUS_LANE modules --------------------------------------------
   -----------------------------------------------------------------------------------------------------------------
   ---------------------------------------------------------
   -----                     Assignements              -----
   ---------------------------------------------------------
   CLK_TX       <= clk_tx_i;
   RST_TXCLK_N  <= rst_sync_gty_n;
   ---------------------------------------------------------
   -----                     Instantiation             -----
   ---------------------------------------------------------
   inst_phy_plus_lane : phy_plus_lane_64b
   port map(
      RST_N                            => RST_N,
      CLK                              => CLK,
      RST_TXCLK_N                      => rst_sync_gty_n,
      LANE_RESET_PPL_OUT               => lane_reset_ppl_out,
      CLK_TX_OUT                       => clk_tx_i,
	   RST_TX_DONE                      => rst_tx_done,
      -- Clock and reset
      ------------------
      CLK_REF_N                        => CLK_REF_N,               -- Clock signal
      CLK_REF_P                        => CLK_REF_P,
      -- FROM Data-link layer
      DATA_TX                          => data_tx_mux,
      CAPABILITY_TX                    => capability_tx_mux,
      NEW_DATA_TX                      => new_data_tx_mux,
      VALID_K_CHARAC_TX                => valid_k_charac_tx_mux,
      FIFO_TX_FULL                     => fifo_tx_full_ppl,
      -- TO Data-link layer
      FIFO_RX_RD_EN                    => fifo_rx_rd_en_demux,
      DATA_RX                          => data_rx_ppl,
      FIFO_RX_EMPTY                    => fifo_rx_empty_ppl,
      FIFO_RX_DATA_VALID               => fifo_rx_data_valid_ppl,
      VALID_K_CHARAC_RX                => valid_k_charac_rx_ppl,
      FAR_END_CAPA_DL                  => far_end_capa_dl_ppl,
      LANE_ACTIVE_DL                   => lane_active_ppl,
      LANE_RESET_DL                    => lane_reset_mux,
      -- FROM/TO Outside
      TX_POS                           => TX_POS,
      TX_NEG                           => TX_NEG,
      RX_POS                           => RX_POS,
      RX_NEG                           => RX_NEG,
      -- PARAMETERS and STATUS
      LANE_START                       => lane_start_ppl,
      AUTOSTART                        => autostart_ppl,
      LANE_RESET                       => lane_reset_ppl,
      PARALLEL_LOOPBACK_EN             => parallel_loopback_en_ppl,
      STANDBY_REASON                   => standby_reason_ppl,
      NEAR_END_SERIAL_LB_EN            => near_end_serial_lb_en_ppl,
      FAR_END_SERIAL_LB_EN             => far_end_serial_lb_en_ppl,
      LANE_STATE                       => lane_state_ppl,
      RX_ERROR_CNT                     => rx_error_cnt_ppl,
      RX_ERROR_OVF                     => rx_error_ovf_ppl,
      LOSS_SIGNAL                      => loss_signal_ppl,
      FAR_END_CAPA                     => far_end_capa_ppl,
      RX_POLARITY                      => rx_polarity_ppl
   );

   inst_mib_phy_plus_lane : mib_phy_plus_lane
   port map(
      -- Parameters From USERAPP/TOP
      LANE_START                       => LANE_START,
      AUTOSTART                        => AUTOSTART,
      LANE_RESET                       => LANE_RESET,
      PARALLEL_LOOPBACK_EN             => PARALLEL_LOOPBACK_EN,
      STANDBY_REASON                   => STANDBY_REASON,
      NEAR_END_SERIAL_LB_EN            => NEAR_END_SERIAL_LB_EN,
      FAR_END_SERIAL_LB_EN             => FAR_END_SERIAL_LB_EN,
      -- Status To USERAPP/TOP
      LANE_STATE                       => LANE_STATE,
      RX_ERROR_CNT                     => RX_ERROR_CNT,
      RX_ERROR_OVF                     => RX_ERROR_OVF,
      LOSS_SIGNAL                      => LOSS_SIGNAL,
      FAR_END_CAPA                     => FAR_END_CAPA,
      RX_POLARITY                      => RX_POLARITY,
      -- Parameters to Module PHY+LANE
      LANE_START_TO_MOD                => lane_start_ppl,
      AUTOSTART_TO_MOD                 => autostart_ppl,
      LANE_RESET_TO_MOD                => lane_reset_ppl,
      PARALLEL_LOOPBACK_EN_TO_MOD      => parallel_loopback_en_ppl,
      STANDBY_REASON_TO_MOD            => standby_reason_ppl,
      NEAR_END_SERIAL_LB_EN_TO_MOD     => near_end_serial_lb_en_ppl,
      FAR_END_SERIAL_LB_EN_TO_MOD      => far_end_serial_lb_en_ppl,
      -- Status from Module PHY+LANE
      LANE_STATE_FROM_MOD              => lane_state_ppl,
      RX_ERROR_CNT_FROM_MOD            => rx_error_cnt_ppl,
      RX_ERROR_OVF_FROM_MOD            => rx_error_ovf_ppl,
      LOSS_SIGNAL_FROM_MOD             => loss_signal_ppl,
      FAR_END_CAPA_FROM_MOD            => far_end_capa_ppl,
      RX_POLARITY_FROM_MOD             => rx_polarity_ppl
   );

end architecture rtl;
