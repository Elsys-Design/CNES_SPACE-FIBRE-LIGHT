// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTHE4_CHANNEL_DEFINES_VH
`else
`define B_GTHE4_CHANNEL_DEFINES_VH

// Look-up table parameters
//

`define GTHE4_CHANNEL_ADDR_N  504
`define GTHE4_CHANNEL_ADDR_SZ 32
`define GTHE4_CHANNEL_DATA_SZ 160

// Attribute addresses
//

`define GTHE4_CHANNEL__ACJTAG_DEBUG_MODE    32'h00000000
`define GTHE4_CHANNEL__ACJTAG_DEBUG_MODE_SZ 1

`define GTHE4_CHANNEL__ACJTAG_MODE    32'h00000001
`define GTHE4_CHANNEL__ACJTAG_MODE_SZ 1

`define GTHE4_CHANNEL__ACJTAG_RESET    32'h00000002
`define GTHE4_CHANNEL__ACJTAG_RESET_SZ 1

`define GTHE4_CHANNEL__ADAPT_CFG0    32'h00000003
`define GTHE4_CHANNEL__ADAPT_CFG0_SZ 16

`define GTHE4_CHANNEL__ADAPT_CFG1    32'h00000004
`define GTHE4_CHANNEL__ADAPT_CFG1_SZ 16

`define GTHE4_CHANNEL__ADAPT_CFG2    32'h00000005
`define GTHE4_CHANNEL__ADAPT_CFG2_SZ 16

`define GTHE4_CHANNEL__ALIGN_COMMA_DOUBLE    32'h00000006
`define GTHE4_CHANNEL__ALIGN_COMMA_DOUBLE_SZ 40

`define GTHE4_CHANNEL__ALIGN_COMMA_ENABLE    32'h00000007
`define GTHE4_CHANNEL__ALIGN_COMMA_ENABLE_SZ 10

`define GTHE4_CHANNEL__ALIGN_COMMA_WORD    32'h00000008
`define GTHE4_CHANNEL__ALIGN_COMMA_WORD_SZ 3

`define GTHE4_CHANNEL__ALIGN_MCOMMA_DET    32'h00000009
`define GTHE4_CHANNEL__ALIGN_MCOMMA_DET_SZ 40

`define GTHE4_CHANNEL__ALIGN_MCOMMA_VALUE    32'h0000000a
`define GTHE4_CHANNEL__ALIGN_MCOMMA_VALUE_SZ 10

`define GTHE4_CHANNEL__ALIGN_PCOMMA_DET    32'h0000000b
`define GTHE4_CHANNEL__ALIGN_PCOMMA_DET_SZ 40

`define GTHE4_CHANNEL__ALIGN_PCOMMA_VALUE    32'h0000000c
`define GTHE4_CHANNEL__ALIGN_PCOMMA_VALUE_SZ 10

`define GTHE4_CHANNEL__A_RXOSCALRESET    32'h0000000d
`define GTHE4_CHANNEL__A_RXOSCALRESET_SZ 1

`define GTHE4_CHANNEL__A_RXPROGDIVRESET    32'h0000000e
`define GTHE4_CHANNEL__A_RXPROGDIVRESET_SZ 1

`define GTHE4_CHANNEL__A_RXTERMINATION    32'h0000000f
`define GTHE4_CHANNEL__A_RXTERMINATION_SZ 1

`define GTHE4_CHANNEL__A_TXDIFFCTRL    32'h00000010
`define GTHE4_CHANNEL__A_TXDIFFCTRL_SZ 5

`define GTHE4_CHANNEL__A_TXPROGDIVRESET    32'h00000011
`define GTHE4_CHANNEL__A_TXPROGDIVRESET_SZ 1

`define GTHE4_CHANNEL__CAPBYPASS_FORCE    32'h00000012
`define GTHE4_CHANNEL__CAPBYPASS_FORCE_SZ 1

`define GTHE4_CHANNEL__CBCC_DATA_SOURCE_SEL    32'h00000013
`define GTHE4_CHANNEL__CBCC_DATA_SOURCE_SEL_SZ 56

`define GTHE4_CHANNEL__CDR_SWAP_MODE_EN    32'h00000014
`define GTHE4_CHANNEL__CDR_SWAP_MODE_EN_SZ 1

`define GTHE4_CHANNEL__CFOK_PWRSVE_EN    32'h00000015
`define GTHE4_CHANNEL__CFOK_PWRSVE_EN_SZ 1

`define GTHE4_CHANNEL__CHAN_BOND_KEEP_ALIGN    32'h00000016
`define GTHE4_CHANNEL__CHAN_BOND_KEEP_ALIGN_SZ 40

`define GTHE4_CHANNEL__CHAN_BOND_MAX_SKEW    32'h00000017
`define GTHE4_CHANNEL__CHAN_BOND_MAX_SKEW_SZ 4

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_1    32'h00000018
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_1_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_2    32'h00000019
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_2_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_3    32'h0000001a
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_3_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_4    32'h0000001b
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_4_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_ENABLE    32'h0000001c
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_1_ENABLE_SZ 4

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_1    32'h0000001d
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_1_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_2    32'h0000001e
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_2_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_3    32'h0000001f
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_3_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_4    32'h00000020
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_4_SZ 10

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_ENABLE    32'h00000021
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_ENABLE_SZ 4

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_USE    32'h00000022
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_2_USE_SZ 40

`define GTHE4_CHANNEL__CHAN_BOND_SEQ_LEN    32'h00000023
`define GTHE4_CHANNEL__CHAN_BOND_SEQ_LEN_SZ 3

`define GTHE4_CHANNEL__CH_HSPMUX    32'h00000024
`define GTHE4_CHANNEL__CH_HSPMUX_SZ 16

`define GTHE4_CHANNEL__CKCAL1_CFG_0    32'h00000025
`define GTHE4_CHANNEL__CKCAL1_CFG_0_SZ 16

`define GTHE4_CHANNEL__CKCAL1_CFG_1    32'h00000026
`define GTHE4_CHANNEL__CKCAL1_CFG_1_SZ 16

`define GTHE4_CHANNEL__CKCAL1_CFG_2    32'h00000027
`define GTHE4_CHANNEL__CKCAL1_CFG_2_SZ 16

`define GTHE4_CHANNEL__CKCAL1_CFG_3    32'h00000028
`define GTHE4_CHANNEL__CKCAL1_CFG_3_SZ 16

`define GTHE4_CHANNEL__CKCAL2_CFG_0    32'h00000029
`define GTHE4_CHANNEL__CKCAL2_CFG_0_SZ 16

`define GTHE4_CHANNEL__CKCAL2_CFG_1    32'h0000002a
`define GTHE4_CHANNEL__CKCAL2_CFG_1_SZ 16

`define GTHE4_CHANNEL__CKCAL2_CFG_2    32'h0000002b
`define GTHE4_CHANNEL__CKCAL2_CFG_2_SZ 16

`define GTHE4_CHANNEL__CKCAL2_CFG_3    32'h0000002c
`define GTHE4_CHANNEL__CKCAL2_CFG_3_SZ 16

`define GTHE4_CHANNEL__CKCAL2_CFG_4    32'h0000002d
`define GTHE4_CHANNEL__CKCAL2_CFG_4_SZ 16

`define GTHE4_CHANNEL__CKCAL_RSVD0    32'h0000002e
`define GTHE4_CHANNEL__CKCAL_RSVD0_SZ 16

`define GTHE4_CHANNEL__CKCAL_RSVD1    32'h0000002f
`define GTHE4_CHANNEL__CKCAL_RSVD1_SZ 16

`define GTHE4_CHANNEL__CLK_CORRECT_USE    32'h00000030
`define GTHE4_CHANNEL__CLK_CORRECT_USE_SZ 40

`define GTHE4_CHANNEL__CLK_COR_KEEP_IDLE    32'h00000031
`define GTHE4_CHANNEL__CLK_COR_KEEP_IDLE_SZ 40

`define GTHE4_CHANNEL__CLK_COR_MAX_LAT    32'h00000032
`define GTHE4_CHANNEL__CLK_COR_MAX_LAT_SZ 6

`define GTHE4_CHANNEL__CLK_COR_MIN_LAT    32'h00000033
`define GTHE4_CHANNEL__CLK_COR_MIN_LAT_SZ 6

`define GTHE4_CHANNEL__CLK_COR_PRECEDENCE    32'h00000034
`define GTHE4_CHANNEL__CLK_COR_PRECEDENCE_SZ 40

`define GTHE4_CHANNEL__CLK_COR_REPEAT_WAIT    32'h00000035
`define GTHE4_CHANNEL__CLK_COR_REPEAT_WAIT_SZ 5

`define GTHE4_CHANNEL__CLK_COR_SEQ_1_1    32'h00000036
`define GTHE4_CHANNEL__CLK_COR_SEQ_1_1_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_1_2    32'h00000037
`define GTHE4_CHANNEL__CLK_COR_SEQ_1_2_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_1_3    32'h00000038
`define GTHE4_CHANNEL__CLK_COR_SEQ_1_3_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_1_4    32'h00000039
`define GTHE4_CHANNEL__CLK_COR_SEQ_1_4_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_1_ENABLE    32'h0000003a
`define GTHE4_CHANNEL__CLK_COR_SEQ_1_ENABLE_SZ 4

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_1    32'h0000003b
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_1_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_2    32'h0000003c
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_2_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_3    32'h0000003d
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_3_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_4    32'h0000003e
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_4_SZ 10

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_ENABLE    32'h0000003f
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_ENABLE_SZ 4

`define GTHE4_CHANNEL__CLK_COR_SEQ_2_USE    32'h00000040
`define GTHE4_CHANNEL__CLK_COR_SEQ_2_USE_SZ 40

`define GTHE4_CHANNEL__CLK_COR_SEQ_LEN    32'h00000041
`define GTHE4_CHANNEL__CLK_COR_SEQ_LEN_SZ 3

`define GTHE4_CHANNEL__CPLL_CFG0    32'h00000042
`define GTHE4_CHANNEL__CPLL_CFG0_SZ 16

`define GTHE4_CHANNEL__CPLL_CFG1    32'h00000043
`define GTHE4_CHANNEL__CPLL_CFG1_SZ 16

`define GTHE4_CHANNEL__CPLL_CFG2    32'h00000044
`define GTHE4_CHANNEL__CPLL_CFG2_SZ 16

`define GTHE4_CHANNEL__CPLL_CFG3    32'h00000045
`define GTHE4_CHANNEL__CPLL_CFG3_SZ 16

`define GTHE4_CHANNEL__CPLL_FBDIV    32'h00000046
`define GTHE4_CHANNEL__CPLL_FBDIV_SZ 5

`define GTHE4_CHANNEL__CPLL_FBDIV_45    32'h00000047
`define GTHE4_CHANNEL__CPLL_FBDIV_45_SZ 3

`define GTHE4_CHANNEL__CPLL_INIT_CFG0    32'h00000048
`define GTHE4_CHANNEL__CPLL_INIT_CFG0_SZ 16

`define GTHE4_CHANNEL__CPLL_LOCK_CFG    32'h00000049
`define GTHE4_CHANNEL__CPLL_LOCK_CFG_SZ 16

`define GTHE4_CHANNEL__CPLL_REFCLK_DIV    32'h0000004a
`define GTHE4_CHANNEL__CPLL_REFCLK_DIV_SZ 5

`define GTHE4_CHANNEL__CTLE3_OCAP_EXT_CTRL    32'h0000004b
`define GTHE4_CHANNEL__CTLE3_OCAP_EXT_CTRL_SZ 3

`define GTHE4_CHANNEL__CTLE3_OCAP_EXT_EN    32'h0000004c
`define GTHE4_CHANNEL__CTLE3_OCAP_EXT_EN_SZ 1

`define GTHE4_CHANNEL__DDI_CTRL    32'h0000004d
`define GTHE4_CHANNEL__DDI_CTRL_SZ 2

`define GTHE4_CHANNEL__DDI_REALIGN_WAIT    32'h0000004e
`define GTHE4_CHANNEL__DDI_REALIGN_WAIT_SZ 5

`define GTHE4_CHANNEL__DEC_MCOMMA_DETECT    32'h0000004f
`define GTHE4_CHANNEL__DEC_MCOMMA_DETECT_SZ 40

`define GTHE4_CHANNEL__DEC_PCOMMA_DETECT    32'h00000050
`define GTHE4_CHANNEL__DEC_PCOMMA_DETECT_SZ 40

`define GTHE4_CHANNEL__DEC_VALID_COMMA_ONLY    32'h00000051
`define GTHE4_CHANNEL__DEC_VALID_COMMA_ONLY_SZ 40

`define GTHE4_CHANNEL__DELAY_ELEC    32'h00000052
`define GTHE4_CHANNEL__DELAY_ELEC_SZ 1

`define GTHE4_CHANNEL__DMONITOR_CFG0    32'h00000053
`define GTHE4_CHANNEL__DMONITOR_CFG0_SZ 10

`define GTHE4_CHANNEL__DMONITOR_CFG1    32'h00000054
`define GTHE4_CHANNEL__DMONITOR_CFG1_SZ 8

`define GTHE4_CHANNEL__ES_CLK_PHASE_SEL    32'h00000055
`define GTHE4_CHANNEL__ES_CLK_PHASE_SEL_SZ 1

`define GTHE4_CHANNEL__ES_CONTROL    32'h00000056
`define GTHE4_CHANNEL__ES_CONTROL_SZ 6

`define GTHE4_CHANNEL__ES_ERRDET_EN    32'h00000057
`define GTHE4_CHANNEL__ES_ERRDET_EN_SZ 40

`define GTHE4_CHANNEL__ES_EYE_SCAN_EN    32'h00000058
`define GTHE4_CHANNEL__ES_EYE_SCAN_EN_SZ 40

`define GTHE4_CHANNEL__ES_HORZ_OFFSET    32'h00000059
`define GTHE4_CHANNEL__ES_HORZ_OFFSET_SZ 12

`define GTHE4_CHANNEL__ES_PRESCALE    32'h0000005a
`define GTHE4_CHANNEL__ES_PRESCALE_SZ 5

`define GTHE4_CHANNEL__ES_QUALIFIER0    32'h0000005b
`define GTHE4_CHANNEL__ES_QUALIFIER0_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER1    32'h0000005c
`define GTHE4_CHANNEL__ES_QUALIFIER1_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER2    32'h0000005d
`define GTHE4_CHANNEL__ES_QUALIFIER2_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER3    32'h0000005e
`define GTHE4_CHANNEL__ES_QUALIFIER3_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER4    32'h0000005f
`define GTHE4_CHANNEL__ES_QUALIFIER4_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER5    32'h00000060
`define GTHE4_CHANNEL__ES_QUALIFIER5_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER6    32'h00000061
`define GTHE4_CHANNEL__ES_QUALIFIER6_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER7    32'h00000062
`define GTHE4_CHANNEL__ES_QUALIFIER7_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER8    32'h00000063
`define GTHE4_CHANNEL__ES_QUALIFIER8_SZ 16

`define GTHE4_CHANNEL__ES_QUALIFIER9    32'h00000064
`define GTHE4_CHANNEL__ES_QUALIFIER9_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK0    32'h00000065
`define GTHE4_CHANNEL__ES_QUAL_MASK0_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK1    32'h00000066
`define GTHE4_CHANNEL__ES_QUAL_MASK1_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK2    32'h00000067
`define GTHE4_CHANNEL__ES_QUAL_MASK2_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK3    32'h00000068
`define GTHE4_CHANNEL__ES_QUAL_MASK3_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK4    32'h00000069
`define GTHE4_CHANNEL__ES_QUAL_MASK4_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK5    32'h0000006a
`define GTHE4_CHANNEL__ES_QUAL_MASK5_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK6    32'h0000006b
`define GTHE4_CHANNEL__ES_QUAL_MASK6_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK7    32'h0000006c
`define GTHE4_CHANNEL__ES_QUAL_MASK7_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK8    32'h0000006d
`define GTHE4_CHANNEL__ES_QUAL_MASK8_SZ 16

`define GTHE4_CHANNEL__ES_QUAL_MASK9    32'h0000006e
`define GTHE4_CHANNEL__ES_QUAL_MASK9_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK0    32'h0000006f
`define GTHE4_CHANNEL__ES_SDATA_MASK0_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK1    32'h00000070
`define GTHE4_CHANNEL__ES_SDATA_MASK1_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK2    32'h00000071
`define GTHE4_CHANNEL__ES_SDATA_MASK2_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK3    32'h00000072
`define GTHE4_CHANNEL__ES_SDATA_MASK3_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK4    32'h00000073
`define GTHE4_CHANNEL__ES_SDATA_MASK4_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK5    32'h00000074
`define GTHE4_CHANNEL__ES_SDATA_MASK5_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK6    32'h00000075
`define GTHE4_CHANNEL__ES_SDATA_MASK6_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK7    32'h00000076
`define GTHE4_CHANNEL__ES_SDATA_MASK7_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK8    32'h00000077
`define GTHE4_CHANNEL__ES_SDATA_MASK8_SZ 16

`define GTHE4_CHANNEL__ES_SDATA_MASK9    32'h00000078
`define GTHE4_CHANNEL__ES_SDATA_MASK9_SZ 16

`define GTHE4_CHANNEL__EYE_SCAN_SWAP_EN    32'h00000079
`define GTHE4_CHANNEL__EYE_SCAN_SWAP_EN_SZ 1

`define GTHE4_CHANNEL__FTS_DESKEW_SEQ_ENABLE    32'h0000007a
`define GTHE4_CHANNEL__FTS_DESKEW_SEQ_ENABLE_SZ 4

`define GTHE4_CHANNEL__FTS_LANE_DESKEW_CFG    32'h0000007b
`define GTHE4_CHANNEL__FTS_LANE_DESKEW_CFG_SZ 4

`define GTHE4_CHANNEL__FTS_LANE_DESKEW_EN    32'h0000007c
`define GTHE4_CHANNEL__FTS_LANE_DESKEW_EN_SZ 40

`define GTHE4_CHANNEL__GEARBOX_MODE    32'h0000007d
`define GTHE4_CHANNEL__GEARBOX_MODE_SZ 5

`define GTHE4_CHANNEL__ISCAN_CK_PH_SEL2    32'h0000007e
`define GTHE4_CHANNEL__ISCAN_CK_PH_SEL2_SZ 1

`define GTHE4_CHANNEL__LOCAL_MASTER    32'h0000007f
`define GTHE4_CHANNEL__LOCAL_MASTER_SZ 1

`define GTHE4_CHANNEL__LPBK_BIAS_CTRL    32'h00000080
`define GTHE4_CHANNEL__LPBK_BIAS_CTRL_SZ 3

`define GTHE4_CHANNEL__LPBK_EN_RCAL_B    32'h00000081
`define GTHE4_CHANNEL__LPBK_EN_RCAL_B_SZ 1

`define GTHE4_CHANNEL__LPBK_EXT_RCAL    32'h00000082
`define GTHE4_CHANNEL__LPBK_EXT_RCAL_SZ 4

`define GTHE4_CHANNEL__LPBK_IND_CTRL0    32'h00000083
`define GTHE4_CHANNEL__LPBK_IND_CTRL0_SZ 3

`define GTHE4_CHANNEL__LPBK_IND_CTRL1    32'h00000084
`define GTHE4_CHANNEL__LPBK_IND_CTRL1_SZ 3

`define GTHE4_CHANNEL__LPBK_IND_CTRL2    32'h00000085
`define GTHE4_CHANNEL__LPBK_IND_CTRL2_SZ 3

`define GTHE4_CHANNEL__LPBK_RG_CTRL    32'h00000086
`define GTHE4_CHANNEL__LPBK_RG_CTRL_SZ 4

`define GTHE4_CHANNEL__OOBDIVCTL    32'h00000087
`define GTHE4_CHANNEL__OOBDIVCTL_SZ 2

`define GTHE4_CHANNEL__OOB_PWRUP    32'h00000088
`define GTHE4_CHANNEL__OOB_PWRUP_SZ 1

`define GTHE4_CHANNEL__PCI3_AUTO_REALIGN    32'h00000089
`define GTHE4_CHANNEL__PCI3_AUTO_REALIGN_SZ 80

`define GTHE4_CHANNEL__PCI3_PIPE_RX_ELECIDLE    32'h0000008a
`define GTHE4_CHANNEL__PCI3_PIPE_RX_ELECIDLE_SZ 1

`define GTHE4_CHANNEL__PCI3_RX_ASYNC_EBUF_BYPASS    32'h0000008b
`define GTHE4_CHANNEL__PCI3_RX_ASYNC_EBUF_BYPASS_SZ 2

`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_EI2_ENABLE    32'h0000008c
`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_EI2_ENABLE_SZ 1

`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_H2L_COUNT    32'h0000008d
`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_H2L_COUNT_SZ 6

`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_H2L_DISABLE    32'h0000008e
`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_H2L_DISABLE_SZ 3

`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_HI_COUNT    32'h0000008f
`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_HI_COUNT_SZ 6

`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_LP4_DISABLE    32'h00000090
`define GTHE4_CHANNEL__PCI3_RX_ELECIDLE_LP4_DISABLE_SZ 1

`define GTHE4_CHANNEL__PCI3_RX_FIFO_DISABLE    32'h00000091
`define GTHE4_CHANNEL__PCI3_RX_FIFO_DISABLE_SZ 1

`define GTHE4_CHANNEL__PCIE3_CLK_COR_EMPTY_THRSH    32'h00000092
`define GTHE4_CHANNEL__PCIE3_CLK_COR_EMPTY_THRSH_SZ 5

`define GTHE4_CHANNEL__PCIE3_CLK_COR_FULL_THRSH    32'h00000093
`define GTHE4_CHANNEL__PCIE3_CLK_COR_FULL_THRSH_SZ 6

`define GTHE4_CHANNEL__PCIE3_CLK_COR_MAX_LAT    32'h00000094
`define GTHE4_CHANNEL__PCIE3_CLK_COR_MAX_LAT_SZ 5

`define GTHE4_CHANNEL__PCIE3_CLK_COR_MIN_LAT    32'h00000095
`define GTHE4_CHANNEL__PCIE3_CLK_COR_MIN_LAT_SZ 5

`define GTHE4_CHANNEL__PCIE3_CLK_COR_THRSH_TIMER    32'h00000096
`define GTHE4_CHANNEL__PCIE3_CLK_COR_THRSH_TIMER_SZ 6

`define GTHE4_CHANNEL__PCIE_BUFG_DIV_CTRL    32'h00000097
`define GTHE4_CHANNEL__PCIE_BUFG_DIV_CTRL_SZ 16

`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN12    32'h00000098
`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN12_SZ 2

`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN3    32'h00000099
`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN3_SZ 2

`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN4    32'h0000009a
`define GTHE4_CHANNEL__PCIE_PLL_SEL_MODE_GEN4_SZ 2

`define GTHE4_CHANNEL__PCIE_RXPCS_CFG_GEN3    32'h0000009b
`define GTHE4_CHANNEL__PCIE_RXPCS_CFG_GEN3_SZ 16

`define GTHE4_CHANNEL__PCIE_RXPMA_CFG    32'h0000009c
`define GTHE4_CHANNEL__PCIE_RXPMA_CFG_SZ 16

`define GTHE4_CHANNEL__PCIE_TXPCS_CFG_GEN3    32'h0000009d
`define GTHE4_CHANNEL__PCIE_TXPCS_CFG_GEN3_SZ 16

`define GTHE4_CHANNEL__PCIE_TXPMA_CFG    32'h0000009e
`define GTHE4_CHANNEL__PCIE_TXPMA_CFG_SZ 16

`define GTHE4_CHANNEL__PCS_PCIE_EN    32'h0000009f
`define GTHE4_CHANNEL__PCS_PCIE_EN_SZ 40

`define GTHE4_CHANNEL__PCS_RSVD0    32'h000000a0
`define GTHE4_CHANNEL__PCS_RSVD0_SZ 16

`define GTHE4_CHANNEL__PD_TRANS_TIME_FROM_P2    32'h000000a1
`define GTHE4_CHANNEL__PD_TRANS_TIME_FROM_P2_SZ 12

`define GTHE4_CHANNEL__PD_TRANS_TIME_NONE_P2    32'h000000a2
`define GTHE4_CHANNEL__PD_TRANS_TIME_NONE_P2_SZ 8

`define GTHE4_CHANNEL__PD_TRANS_TIME_TO_P2    32'h000000a3
`define GTHE4_CHANNEL__PD_TRANS_TIME_TO_P2_SZ 8

`define GTHE4_CHANNEL__PREIQ_FREQ_BST    32'h000000a4
`define GTHE4_CHANNEL__PREIQ_FREQ_BST_SZ 2

`define GTHE4_CHANNEL__PROCESS_PAR    32'h000000a5
`define GTHE4_CHANNEL__PROCESS_PAR_SZ 3

`define GTHE4_CHANNEL__RATE_SW_USE_DRP    32'h000000a6
`define GTHE4_CHANNEL__RATE_SW_USE_DRP_SZ 1

`define GTHE4_CHANNEL__RCLK_SIPO_DLY_ENB    32'h000000a7
`define GTHE4_CHANNEL__RCLK_SIPO_DLY_ENB_SZ 1

`define GTHE4_CHANNEL__RCLK_SIPO_INV_EN    32'h000000a8
`define GTHE4_CHANNEL__RCLK_SIPO_INV_EN_SZ 1

`define GTHE4_CHANNEL__RESET_POWERSAVE_DISABLE    32'h000000a9
`define GTHE4_CHANNEL__RESET_POWERSAVE_DISABLE_SZ 1

`define GTHE4_CHANNEL__RTX_BUF_CML_CTRL    32'h000000aa
`define GTHE4_CHANNEL__RTX_BUF_CML_CTRL_SZ 3

`define GTHE4_CHANNEL__RTX_BUF_TERM_CTRL    32'h000000ab
`define GTHE4_CHANNEL__RTX_BUF_TERM_CTRL_SZ 2

`define GTHE4_CHANNEL__RXBUFRESET_TIME    32'h000000ac
`define GTHE4_CHANNEL__RXBUFRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXBUF_ADDR_MODE    32'h000000ad
`define GTHE4_CHANNEL__RXBUF_ADDR_MODE_SZ 32

`define GTHE4_CHANNEL__RXBUF_EIDLE_HI_CNT    32'h000000ae
`define GTHE4_CHANNEL__RXBUF_EIDLE_HI_CNT_SZ 4

`define GTHE4_CHANNEL__RXBUF_EIDLE_LO_CNT    32'h000000af
`define GTHE4_CHANNEL__RXBUF_EIDLE_LO_CNT_SZ 4

`define GTHE4_CHANNEL__RXBUF_EN    32'h000000b0
`define GTHE4_CHANNEL__RXBUF_EN_SZ 40

`define GTHE4_CHANNEL__RXBUF_RESET_ON_CB_CHANGE    32'h000000b1
`define GTHE4_CHANNEL__RXBUF_RESET_ON_CB_CHANGE_SZ 40

`define GTHE4_CHANNEL__RXBUF_RESET_ON_COMMAALIGN    32'h000000b2
`define GTHE4_CHANNEL__RXBUF_RESET_ON_COMMAALIGN_SZ 40

`define GTHE4_CHANNEL__RXBUF_RESET_ON_EIDLE    32'h000000b3
`define GTHE4_CHANNEL__RXBUF_RESET_ON_EIDLE_SZ 40

`define GTHE4_CHANNEL__RXBUF_RESET_ON_RATE_CHANGE    32'h000000b4
`define GTHE4_CHANNEL__RXBUF_RESET_ON_RATE_CHANGE_SZ 40

`define GTHE4_CHANNEL__RXBUF_THRESH_OVFLW    32'h000000b5
`define GTHE4_CHANNEL__RXBUF_THRESH_OVFLW_SZ 6

`define GTHE4_CHANNEL__RXBUF_THRESH_OVRD    32'h000000b6
`define GTHE4_CHANNEL__RXBUF_THRESH_OVRD_SZ 40

`define GTHE4_CHANNEL__RXBUF_THRESH_UNDFLW    32'h000000b7
`define GTHE4_CHANNEL__RXBUF_THRESH_UNDFLW_SZ 6

`define GTHE4_CHANNEL__RXCDRFREQRESET_TIME    32'h000000b8
`define GTHE4_CHANNEL__RXCDRFREQRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXCDRPHRESET_TIME    32'h000000b9
`define GTHE4_CHANNEL__RXCDRPHRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXCDR_CFG0    32'h000000ba
`define GTHE4_CHANNEL__RXCDR_CFG0_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG0_GEN3    32'h000000bb
`define GTHE4_CHANNEL__RXCDR_CFG0_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG1    32'h000000bc
`define GTHE4_CHANNEL__RXCDR_CFG1_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG1_GEN3    32'h000000bd
`define GTHE4_CHANNEL__RXCDR_CFG1_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG2    32'h000000be
`define GTHE4_CHANNEL__RXCDR_CFG2_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG2_GEN2    32'h000000bf
`define GTHE4_CHANNEL__RXCDR_CFG2_GEN2_SZ 10

`define GTHE4_CHANNEL__RXCDR_CFG2_GEN3    32'h000000c0
`define GTHE4_CHANNEL__RXCDR_CFG2_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG2_GEN4    32'h000000c1
`define GTHE4_CHANNEL__RXCDR_CFG2_GEN4_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG3    32'h000000c2
`define GTHE4_CHANNEL__RXCDR_CFG3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG3_GEN2    32'h000000c3
`define GTHE4_CHANNEL__RXCDR_CFG3_GEN2_SZ 6

`define GTHE4_CHANNEL__RXCDR_CFG3_GEN3    32'h000000c4
`define GTHE4_CHANNEL__RXCDR_CFG3_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG3_GEN4    32'h000000c5
`define GTHE4_CHANNEL__RXCDR_CFG3_GEN4_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG4    32'h000000c6
`define GTHE4_CHANNEL__RXCDR_CFG4_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG4_GEN3    32'h000000c7
`define GTHE4_CHANNEL__RXCDR_CFG4_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG5    32'h000000c8
`define GTHE4_CHANNEL__RXCDR_CFG5_SZ 16

`define GTHE4_CHANNEL__RXCDR_CFG5_GEN3    32'h000000c9
`define GTHE4_CHANNEL__RXCDR_CFG5_GEN3_SZ 16

`define GTHE4_CHANNEL__RXCDR_FR_RESET_ON_EIDLE    32'h000000ca
`define GTHE4_CHANNEL__RXCDR_FR_RESET_ON_EIDLE_SZ 1

`define GTHE4_CHANNEL__RXCDR_HOLD_DURING_EIDLE    32'h000000cb
`define GTHE4_CHANNEL__RXCDR_HOLD_DURING_EIDLE_SZ 1

`define GTHE4_CHANNEL__RXCDR_LOCK_CFG0    32'h000000cc
`define GTHE4_CHANNEL__RXCDR_LOCK_CFG0_SZ 16

`define GTHE4_CHANNEL__RXCDR_LOCK_CFG1    32'h000000cd
`define GTHE4_CHANNEL__RXCDR_LOCK_CFG1_SZ 16

`define GTHE4_CHANNEL__RXCDR_LOCK_CFG2    32'h000000ce
`define GTHE4_CHANNEL__RXCDR_LOCK_CFG2_SZ 16

`define GTHE4_CHANNEL__RXCDR_LOCK_CFG3    32'h000000cf
`define GTHE4_CHANNEL__RXCDR_LOCK_CFG3_SZ 16

`define GTHE4_CHANNEL__RXCDR_LOCK_CFG4    32'h000000d0
`define GTHE4_CHANNEL__RXCDR_LOCK_CFG4_SZ 16

`define GTHE4_CHANNEL__RXCDR_PH_RESET_ON_EIDLE    32'h000000d1
`define GTHE4_CHANNEL__RXCDR_PH_RESET_ON_EIDLE_SZ 1

`define GTHE4_CHANNEL__RXCFOK_CFG0    32'h000000d2
`define GTHE4_CHANNEL__RXCFOK_CFG0_SZ 16

`define GTHE4_CHANNEL__RXCFOK_CFG1    32'h000000d3
`define GTHE4_CHANNEL__RXCFOK_CFG1_SZ 16

`define GTHE4_CHANNEL__RXCFOK_CFG2    32'h000000d4
`define GTHE4_CHANNEL__RXCFOK_CFG2_SZ 16

`define GTHE4_CHANNEL__RXCKCAL1_IQ_LOOP_RST_CFG    32'h000000d5
`define GTHE4_CHANNEL__RXCKCAL1_IQ_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL1_I_LOOP_RST_CFG    32'h000000d6
`define GTHE4_CHANNEL__RXCKCAL1_I_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL1_Q_LOOP_RST_CFG    32'h000000d7
`define GTHE4_CHANNEL__RXCKCAL1_Q_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL2_DX_LOOP_RST_CFG    32'h000000d8
`define GTHE4_CHANNEL__RXCKCAL2_DX_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL2_D_LOOP_RST_CFG    32'h000000d9
`define GTHE4_CHANNEL__RXCKCAL2_D_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL2_S_LOOP_RST_CFG    32'h000000da
`define GTHE4_CHANNEL__RXCKCAL2_S_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXCKCAL2_X_LOOP_RST_CFG    32'h000000db
`define GTHE4_CHANNEL__RXCKCAL2_X_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__RXDFELPMRESET_TIME    32'h000000dc
`define GTHE4_CHANNEL__RXDFELPMRESET_TIME_SZ 7

`define GTHE4_CHANNEL__RXDFELPM_KL_CFG0    32'h000000dd
`define GTHE4_CHANNEL__RXDFELPM_KL_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFELPM_KL_CFG1    32'h000000de
`define GTHE4_CHANNEL__RXDFELPM_KL_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFELPM_KL_CFG2    32'h000000df
`define GTHE4_CHANNEL__RXDFELPM_KL_CFG2_SZ 16

`define GTHE4_CHANNEL__RXDFE_CFG0    32'h000000e0
`define GTHE4_CHANNEL__RXDFE_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_CFG1    32'h000000e1
`define GTHE4_CHANNEL__RXDFE_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_GC_CFG0    32'h000000e2
`define GTHE4_CHANNEL__RXDFE_GC_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_GC_CFG1    32'h000000e3
`define GTHE4_CHANNEL__RXDFE_GC_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_GC_CFG2    32'h000000e4
`define GTHE4_CHANNEL__RXDFE_GC_CFG2_SZ 16

`define GTHE4_CHANNEL__RXDFE_H2_CFG0    32'h000000e5
`define GTHE4_CHANNEL__RXDFE_H2_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H2_CFG1    32'h000000e6
`define GTHE4_CHANNEL__RXDFE_H2_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H3_CFG0    32'h000000e7
`define GTHE4_CHANNEL__RXDFE_H3_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H3_CFG1    32'h000000e8
`define GTHE4_CHANNEL__RXDFE_H3_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H4_CFG0    32'h000000e9
`define GTHE4_CHANNEL__RXDFE_H4_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H4_CFG1    32'h000000ea
`define GTHE4_CHANNEL__RXDFE_H4_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H5_CFG0    32'h000000eb
`define GTHE4_CHANNEL__RXDFE_H5_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H5_CFG1    32'h000000ec
`define GTHE4_CHANNEL__RXDFE_H5_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H6_CFG0    32'h000000ed
`define GTHE4_CHANNEL__RXDFE_H6_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H6_CFG1    32'h000000ee
`define GTHE4_CHANNEL__RXDFE_H6_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H7_CFG0    32'h000000ef
`define GTHE4_CHANNEL__RXDFE_H7_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H7_CFG1    32'h000000f0
`define GTHE4_CHANNEL__RXDFE_H7_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H8_CFG0    32'h000000f1
`define GTHE4_CHANNEL__RXDFE_H8_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H8_CFG1    32'h000000f2
`define GTHE4_CHANNEL__RXDFE_H8_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_H9_CFG0    32'h000000f3
`define GTHE4_CHANNEL__RXDFE_H9_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_H9_CFG1    32'h000000f4
`define GTHE4_CHANNEL__RXDFE_H9_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HA_CFG0    32'h000000f5
`define GTHE4_CHANNEL__RXDFE_HA_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HA_CFG1    32'h000000f6
`define GTHE4_CHANNEL__RXDFE_HA_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HB_CFG0    32'h000000f7
`define GTHE4_CHANNEL__RXDFE_HB_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HB_CFG1    32'h000000f8
`define GTHE4_CHANNEL__RXDFE_HB_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HC_CFG0    32'h000000f9
`define GTHE4_CHANNEL__RXDFE_HC_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HC_CFG1    32'h000000fa
`define GTHE4_CHANNEL__RXDFE_HC_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HD_CFG0    32'h000000fb
`define GTHE4_CHANNEL__RXDFE_HD_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HD_CFG1    32'h000000fc
`define GTHE4_CHANNEL__RXDFE_HD_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HE_CFG0    32'h000000fd
`define GTHE4_CHANNEL__RXDFE_HE_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HE_CFG1    32'h000000fe
`define GTHE4_CHANNEL__RXDFE_HE_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_HF_CFG0    32'h000000ff
`define GTHE4_CHANNEL__RXDFE_HF_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_HF_CFG1    32'h00000100
`define GTHE4_CHANNEL__RXDFE_HF_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_KH_CFG0    32'h00000101
`define GTHE4_CHANNEL__RXDFE_KH_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_KH_CFG1    32'h00000102
`define GTHE4_CHANNEL__RXDFE_KH_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_KH_CFG2    32'h00000103
`define GTHE4_CHANNEL__RXDFE_KH_CFG2_SZ 16

`define GTHE4_CHANNEL__RXDFE_KH_CFG3    32'h00000104
`define GTHE4_CHANNEL__RXDFE_KH_CFG3_SZ 16

`define GTHE4_CHANNEL__RXDFE_OS_CFG0    32'h00000105
`define GTHE4_CHANNEL__RXDFE_OS_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_OS_CFG1    32'h00000106
`define GTHE4_CHANNEL__RXDFE_OS_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_PWR_SAVING    32'h00000107
`define GTHE4_CHANNEL__RXDFE_PWR_SAVING_SZ 1

`define GTHE4_CHANNEL__RXDFE_UT_CFG0    32'h00000108
`define GTHE4_CHANNEL__RXDFE_UT_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_UT_CFG1    32'h00000109
`define GTHE4_CHANNEL__RXDFE_UT_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDFE_UT_CFG2    32'h0000010a
`define GTHE4_CHANNEL__RXDFE_UT_CFG2_SZ 16

`define GTHE4_CHANNEL__RXDFE_VP_CFG0    32'h0000010b
`define GTHE4_CHANNEL__RXDFE_VP_CFG0_SZ 16

`define GTHE4_CHANNEL__RXDFE_VP_CFG1    32'h0000010c
`define GTHE4_CHANNEL__RXDFE_VP_CFG1_SZ 16

`define GTHE4_CHANNEL__RXDLY_CFG    32'h0000010d
`define GTHE4_CHANNEL__RXDLY_CFG_SZ 16

`define GTHE4_CHANNEL__RXDLY_LCFG    32'h0000010e
`define GTHE4_CHANNEL__RXDLY_LCFG_SZ 16

`define GTHE4_CHANNEL__RXELECIDLE_CFG    32'h0000010f
`define GTHE4_CHANNEL__RXELECIDLE_CFG_SZ 72

`define GTHE4_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR    32'h00000110
`define GTHE4_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR_SZ 3

`define GTHE4_CHANNEL__RXGEARBOX_EN    32'h00000111
`define GTHE4_CHANNEL__RXGEARBOX_EN_SZ 40

`define GTHE4_CHANNEL__RXISCANRESET_TIME    32'h00000112
`define GTHE4_CHANNEL__RXISCANRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXLPM_CFG    32'h00000113
`define GTHE4_CHANNEL__RXLPM_CFG_SZ 16

`define GTHE4_CHANNEL__RXLPM_GC_CFG    32'h00000114
`define GTHE4_CHANNEL__RXLPM_GC_CFG_SZ 16

`define GTHE4_CHANNEL__RXLPM_KH_CFG0    32'h00000115
`define GTHE4_CHANNEL__RXLPM_KH_CFG0_SZ 16

`define GTHE4_CHANNEL__RXLPM_KH_CFG1    32'h00000116
`define GTHE4_CHANNEL__RXLPM_KH_CFG1_SZ 16

`define GTHE4_CHANNEL__RXLPM_OS_CFG0    32'h00000117
`define GTHE4_CHANNEL__RXLPM_OS_CFG0_SZ 16

`define GTHE4_CHANNEL__RXLPM_OS_CFG1    32'h00000118
`define GTHE4_CHANNEL__RXLPM_OS_CFG1_SZ 16

`define GTHE4_CHANNEL__RXOOB_CFG    32'h00000119
`define GTHE4_CHANNEL__RXOOB_CFG_SZ 9

`define GTHE4_CHANNEL__RXOOB_CLK_CFG    32'h0000011a
`define GTHE4_CHANNEL__RXOOB_CLK_CFG_SZ 48

`define GTHE4_CHANNEL__RXOSCALRESET_TIME    32'h0000011b
`define GTHE4_CHANNEL__RXOSCALRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXOUT_DIV    32'h0000011c
`define GTHE4_CHANNEL__RXOUT_DIV_SZ 5

`define GTHE4_CHANNEL__RXPCSRESET_TIME    32'h0000011d
`define GTHE4_CHANNEL__RXPCSRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXPHBEACON_CFG    32'h0000011e
`define GTHE4_CHANNEL__RXPHBEACON_CFG_SZ 16

`define GTHE4_CHANNEL__RXPHDLY_CFG    32'h0000011f
`define GTHE4_CHANNEL__RXPHDLY_CFG_SZ 16

`define GTHE4_CHANNEL__RXPHSAMP_CFG    32'h00000120
`define GTHE4_CHANNEL__RXPHSAMP_CFG_SZ 16

`define GTHE4_CHANNEL__RXPHSLIP_CFG    32'h00000121
`define GTHE4_CHANNEL__RXPHSLIP_CFG_SZ 16

`define GTHE4_CHANNEL__RXPH_MONITOR_SEL    32'h00000122
`define GTHE4_CHANNEL__RXPH_MONITOR_SEL_SZ 5

`define GTHE4_CHANNEL__RXPI_AUTO_BW_SEL_BYPASS    32'h00000123
`define GTHE4_CHANNEL__RXPI_AUTO_BW_SEL_BYPASS_SZ 1

`define GTHE4_CHANNEL__RXPI_CFG0    32'h00000124
`define GTHE4_CHANNEL__RXPI_CFG0_SZ 16

`define GTHE4_CHANNEL__RXPI_CFG1    32'h00000125
`define GTHE4_CHANNEL__RXPI_CFG1_SZ 16

`define GTHE4_CHANNEL__RXPI_LPM    32'h00000126
`define GTHE4_CHANNEL__RXPI_LPM_SZ 1

`define GTHE4_CHANNEL__RXPI_SEL_LC    32'h00000127
`define GTHE4_CHANNEL__RXPI_SEL_LC_SZ 2

`define GTHE4_CHANNEL__RXPI_STARTCODE    32'h00000128
`define GTHE4_CHANNEL__RXPI_STARTCODE_SZ 2

`define GTHE4_CHANNEL__RXPI_VREFSEL    32'h00000129
`define GTHE4_CHANNEL__RXPI_VREFSEL_SZ 1

`define GTHE4_CHANNEL__RXPMACLK_SEL    32'h0000012a
`define GTHE4_CHANNEL__RXPMACLK_SEL_SZ 64

`define GTHE4_CHANNEL__RXPMARESET_TIME    32'h0000012b
`define GTHE4_CHANNEL__RXPMARESET_TIME_SZ 5

`define GTHE4_CHANNEL__RXPRBS_ERR_LOOPBACK    32'h0000012c
`define GTHE4_CHANNEL__RXPRBS_ERR_LOOPBACK_SZ 1

`define GTHE4_CHANNEL__RXPRBS_LINKACQ_CNT    32'h0000012d
`define GTHE4_CHANNEL__RXPRBS_LINKACQ_CNT_SZ 8

`define GTHE4_CHANNEL__RXREFCLKDIV2_SEL    32'h0000012e
`define GTHE4_CHANNEL__RXREFCLKDIV2_SEL_SZ 1

`define GTHE4_CHANNEL__RXSLIDE_AUTO_WAIT    32'h0000012f
`define GTHE4_CHANNEL__RXSLIDE_AUTO_WAIT_SZ 4

`define GTHE4_CHANNEL__RXSLIDE_MODE    32'h00000130
`define GTHE4_CHANNEL__RXSLIDE_MODE_SZ 32

`define GTHE4_CHANNEL__RXSYNC_MULTILANE    32'h00000131
`define GTHE4_CHANNEL__RXSYNC_MULTILANE_SZ 1

`define GTHE4_CHANNEL__RXSYNC_OVRD    32'h00000132
`define GTHE4_CHANNEL__RXSYNC_OVRD_SZ 1

`define GTHE4_CHANNEL__RXSYNC_SKIP_DA    32'h00000133
`define GTHE4_CHANNEL__RXSYNC_SKIP_DA_SZ 1

`define GTHE4_CHANNEL__RX_AFE_CM_EN    32'h00000134
`define GTHE4_CHANNEL__RX_AFE_CM_EN_SZ 1

`define GTHE4_CHANNEL__RX_BIAS_CFG0    32'h00000135
`define GTHE4_CHANNEL__RX_BIAS_CFG0_SZ 16

`define GTHE4_CHANNEL__RX_BUFFER_CFG    32'h00000136
`define GTHE4_CHANNEL__RX_BUFFER_CFG_SZ 6

`define GTHE4_CHANNEL__RX_CAPFF_SARC_ENB    32'h00000137
`define GTHE4_CHANNEL__RX_CAPFF_SARC_ENB_SZ 1

`define GTHE4_CHANNEL__RX_CLK25_DIV    32'h00000138
`define GTHE4_CHANNEL__RX_CLK25_DIV_SZ 6

`define GTHE4_CHANNEL__RX_CLKMUX_EN    32'h00000139
`define GTHE4_CHANNEL__RX_CLKMUX_EN_SZ 1

`define GTHE4_CHANNEL__RX_CLK_SLIP_OVRD    32'h0000013a
`define GTHE4_CHANNEL__RX_CLK_SLIP_OVRD_SZ 5

`define GTHE4_CHANNEL__RX_CM_BUF_CFG    32'h0000013b
`define GTHE4_CHANNEL__RX_CM_BUF_CFG_SZ 4

`define GTHE4_CHANNEL__RX_CM_BUF_PD    32'h0000013c
`define GTHE4_CHANNEL__RX_CM_BUF_PD_SZ 1

`define GTHE4_CHANNEL__RX_CM_SEL    32'h0000013d
`define GTHE4_CHANNEL__RX_CM_SEL_SZ 2

`define GTHE4_CHANNEL__RX_CM_TRIM    32'h0000013e
`define GTHE4_CHANNEL__RX_CM_TRIM_SZ 4

`define GTHE4_CHANNEL__RX_CTLE3_LPF    32'h0000013f
`define GTHE4_CHANNEL__RX_CTLE3_LPF_SZ 8

`define GTHE4_CHANNEL__RX_DATA_WIDTH    32'h00000140
`define GTHE4_CHANNEL__RX_DATA_WIDTH_SZ 8

`define GTHE4_CHANNEL__RX_DDI_SEL    32'h00000141
`define GTHE4_CHANNEL__RX_DDI_SEL_SZ 6

`define GTHE4_CHANNEL__RX_DEFER_RESET_BUF_EN    32'h00000142
`define GTHE4_CHANNEL__RX_DEFER_RESET_BUF_EN_SZ 40

`define GTHE4_CHANNEL__RX_DEGEN_CTRL    32'h00000143
`define GTHE4_CHANNEL__RX_DEGEN_CTRL_SZ 3

`define GTHE4_CHANNEL__RX_DFELPM_CFG0    32'h00000144
`define GTHE4_CHANNEL__RX_DFELPM_CFG0_SZ 4

`define GTHE4_CHANNEL__RX_DFELPM_CFG1    32'h00000145
`define GTHE4_CHANNEL__RX_DFELPM_CFG1_SZ 1

`define GTHE4_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN    32'h00000146
`define GTHE4_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN_SZ 1

`define GTHE4_CHANNEL__RX_DFE_AGC_CFG0    32'h00000147
`define GTHE4_CHANNEL__RX_DFE_AGC_CFG0_SZ 2

`define GTHE4_CHANNEL__RX_DFE_AGC_CFG1    32'h00000148
`define GTHE4_CHANNEL__RX_DFE_AGC_CFG1_SZ 3

`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KH_CFG0    32'h00000149
`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KH_CFG0_SZ 2

`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KH_CFG1    32'h0000014a
`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KH_CFG1_SZ 3

`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KL_CFG0    32'h0000014b
`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KL_CFG0_SZ 2

`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KL_CFG1    32'h0000014c
`define GTHE4_CHANNEL__RX_DFE_KL_LPM_KL_CFG1_SZ 3

`define GTHE4_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE    32'h0000014d
`define GTHE4_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE_SZ 1

`define GTHE4_CHANNEL__RX_DISPERR_SEQ_MATCH    32'h0000014e
`define GTHE4_CHANNEL__RX_DISPERR_SEQ_MATCH_SZ 40

`define GTHE4_CHANNEL__RX_DIV2_MODE_B    32'h0000014f
`define GTHE4_CHANNEL__RX_DIV2_MODE_B_SZ 1

`define GTHE4_CHANNEL__RX_DIVRESET_TIME    32'h00000150
`define GTHE4_CHANNEL__RX_DIVRESET_TIME_SZ 5

`define GTHE4_CHANNEL__RX_EN_CTLE_RCAL_B    32'h00000151
`define GTHE4_CHANNEL__RX_EN_CTLE_RCAL_B_SZ 1

`define GTHE4_CHANNEL__RX_EN_HI_LR    32'h00000152
`define GTHE4_CHANNEL__RX_EN_HI_LR_SZ 1

`define GTHE4_CHANNEL__RX_EXT_RL_CTRL    32'h00000153
`define GTHE4_CHANNEL__RX_EXT_RL_CTRL_SZ 9

`define GTHE4_CHANNEL__RX_EYESCAN_VS_CODE    32'h00000154
`define GTHE4_CHANNEL__RX_EYESCAN_VS_CODE_SZ 7

`define GTHE4_CHANNEL__RX_EYESCAN_VS_NEG_DIR    32'h00000155
`define GTHE4_CHANNEL__RX_EYESCAN_VS_NEG_DIR_SZ 1

`define GTHE4_CHANNEL__RX_EYESCAN_VS_RANGE    32'h00000156
`define GTHE4_CHANNEL__RX_EYESCAN_VS_RANGE_SZ 2

`define GTHE4_CHANNEL__RX_EYESCAN_VS_UT_SIGN    32'h00000157
`define GTHE4_CHANNEL__RX_EYESCAN_VS_UT_SIGN_SZ 1

`define GTHE4_CHANNEL__RX_FABINT_USRCLK_FLOP    32'h00000158
`define GTHE4_CHANNEL__RX_FABINT_USRCLK_FLOP_SZ 1

`define GTHE4_CHANNEL__RX_INT_DATAWIDTH    32'h00000159
`define GTHE4_CHANNEL__RX_INT_DATAWIDTH_SZ 2

`define GTHE4_CHANNEL__RX_PMA_POWER_SAVE    32'h0000015a
`define GTHE4_CHANNEL__RX_PMA_POWER_SAVE_SZ 1

`define GTHE4_CHANNEL__RX_PMA_RSV0    32'h0000015b
`define GTHE4_CHANNEL__RX_PMA_RSV0_SZ 16

`define GTHE4_CHANNEL__RX_PROGDIV_CFG    32'h0000015c
`define GTHE4_CHANNEL__RX_PROGDIV_CFG_SZ 64

`define GTHE4_CHANNEL__RX_PROGDIV_RATE    32'h0000015d
`define GTHE4_CHANNEL__RX_PROGDIV_RATE_SZ 16

`define GTHE4_CHANNEL__RX_RESLOAD_CTRL    32'h0000015e
`define GTHE4_CHANNEL__RX_RESLOAD_CTRL_SZ 4

`define GTHE4_CHANNEL__RX_RESLOAD_OVRD    32'h0000015f
`define GTHE4_CHANNEL__RX_RESLOAD_OVRD_SZ 1

`define GTHE4_CHANNEL__RX_SAMPLE_PERIOD    32'h00000160
`define GTHE4_CHANNEL__RX_SAMPLE_PERIOD_SZ 3

`define GTHE4_CHANNEL__RX_SIG_VALID_DLY    32'h00000161
`define GTHE4_CHANNEL__RX_SIG_VALID_DLY_SZ 6

`define GTHE4_CHANNEL__RX_SUM_DFETAPREP_EN    32'h00000162
`define GTHE4_CHANNEL__RX_SUM_DFETAPREP_EN_SZ 1

`define GTHE4_CHANNEL__RX_SUM_IREF_TUNE    32'h00000163
`define GTHE4_CHANNEL__RX_SUM_IREF_TUNE_SZ 4

`define GTHE4_CHANNEL__RX_SUM_RESLOAD_CTRL    32'h00000164
`define GTHE4_CHANNEL__RX_SUM_RESLOAD_CTRL_SZ 4

`define GTHE4_CHANNEL__RX_SUM_VCMTUNE    32'h00000165
`define GTHE4_CHANNEL__RX_SUM_VCMTUNE_SZ 4

`define GTHE4_CHANNEL__RX_SUM_VCM_OVWR    32'h00000166
`define GTHE4_CHANNEL__RX_SUM_VCM_OVWR_SZ 1

`define GTHE4_CHANNEL__RX_SUM_VREF_TUNE    32'h00000167
`define GTHE4_CHANNEL__RX_SUM_VREF_TUNE_SZ 3

`define GTHE4_CHANNEL__RX_TUNE_AFE_OS    32'h00000168
`define GTHE4_CHANNEL__RX_TUNE_AFE_OS_SZ 2

`define GTHE4_CHANNEL__RX_VREG_CTRL    32'h00000169
`define GTHE4_CHANNEL__RX_VREG_CTRL_SZ 3

`define GTHE4_CHANNEL__RX_VREG_PDB    32'h0000016a
`define GTHE4_CHANNEL__RX_VREG_PDB_SZ 1

`define GTHE4_CHANNEL__RX_WIDEMODE_CDR    32'h0000016b
`define GTHE4_CHANNEL__RX_WIDEMODE_CDR_SZ 2

`define GTHE4_CHANNEL__RX_WIDEMODE_CDR_GEN3    32'h0000016c
`define GTHE4_CHANNEL__RX_WIDEMODE_CDR_GEN3_SZ 2

`define GTHE4_CHANNEL__RX_WIDEMODE_CDR_GEN4    32'h0000016d
`define GTHE4_CHANNEL__RX_WIDEMODE_CDR_GEN4_SZ 2

`define GTHE4_CHANNEL__RX_XCLK_SEL    32'h0000016e
`define GTHE4_CHANNEL__RX_XCLK_SEL_SZ 40

`define GTHE4_CHANNEL__RX_XMODE_SEL    32'h0000016f
`define GTHE4_CHANNEL__RX_XMODE_SEL_SZ 1

`define GTHE4_CHANNEL__SAMPLE_CLK_PHASE    32'h00000170
`define GTHE4_CHANNEL__SAMPLE_CLK_PHASE_SZ 1

`define GTHE4_CHANNEL__SAS_12G_MODE    32'h00000171
`define GTHE4_CHANNEL__SAS_12G_MODE_SZ 1

`define GTHE4_CHANNEL__SATA_BURST_SEQ_LEN    32'h00000172
`define GTHE4_CHANNEL__SATA_BURST_SEQ_LEN_SZ 4

`define GTHE4_CHANNEL__SATA_BURST_VAL    32'h00000173
`define GTHE4_CHANNEL__SATA_BURST_VAL_SZ 3

`define GTHE4_CHANNEL__SATA_CPLL_CFG    32'h00000174
`define GTHE4_CHANNEL__SATA_CPLL_CFG_SZ 88

`define GTHE4_CHANNEL__SATA_EIDLE_VAL    32'h00000175
`define GTHE4_CHANNEL__SATA_EIDLE_VAL_SZ 3

`define GTHE4_CHANNEL__SHOW_REALIGN_COMMA    32'h00000176
`define GTHE4_CHANNEL__SHOW_REALIGN_COMMA_SZ 40

`define GTHE4_CHANNEL__SIM_DEVICE    32'h00000177
`define GTHE4_CHANNEL__SIM_DEVICE_SZ 160

`define GTHE4_CHANNEL__SIM_MODE    32'h00000178
`define GTHE4_CHANNEL__SIM_MODE_SZ 48

`define GTHE4_CHANNEL__SIM_RECEIVER_DETECT_PASS    32'h00000179
`define GTHE4_CHANNEL__SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTHE4_CHANNEL__SIM_RESET_SPEEDUP    32'h0000017a
`define GTHE4_CHANNEL__SIM_RESET_SPEEDUP_SZ 40

`define GTHE4_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL    32'h0000017b
`define GTHE4_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTHE4_CHANNEL__SRSTMODE    32'h0000017c
`define GTHE4_CHANNEL__SRSTMODE_SZ 1

`define GTHE4_CHANNEL__TAPDLY_SET_TX    32'h0000017d
`define GTHE4_CHANNEL__TAPDLY_SET_TX_SZ 2

`define GTHE4_CHANNEL__TEMPERATURE_PAR    32'h0000017e
`define GTHE4_CHANNEL__TEMPERATURE_PAR_SZ 4

`define GTHE4_CHANNEL__TERM_RCAL_CFG    32'h0000017f
`define GTHE4_CHANNEL__TERM_RCAL_CFG_SZ 15

`define GTHE4_CHANNEL__TERM_RCAL_OVRD    32'h00000180
`define GTHE4_CHANNEL__TERM_RCAL_OVRD_SZ 3

`define GTHE4_CHANNEL__TRANS_TIME_RATE    32'h00000181
`define GTHE4_CHANNEL__TRANS_TIME_RATE_SZ 8

`define GTHE4_CHANNEL__TST_RSV0    32'h00000182
`define GTHE4_CHANNEL__TST_RSV0_SZ 8

`define GTHE4_CHANNEL__TST_RSV1    32'h00000183
`define GTHE4_CHANNEL__TST_RSV1_SZ 8

`define GTHE4_CHANNEL__TXBUF_EN    32'h00000184
`define GTHE4_CHANNEL__TXBUF_EN_SZ 40

`define GTHE4_CHANNEL__TXBUF_RESET_ON_RATE_CHANGE    32'h00000185
`define GTHE4_CHANNEL__TXBUF_RESET_ON_RATE_CHANGE_SZ 40

`define GTHE4_CHANNEL__TXDLY_CFG    32'h00000186
`define GTHE4_CHANNEL__TXDLY_CFG_SZ 16

`define GTHE4_CHANNEL__TXDLY_LCFG    32'h00000187
`define GTHE4_CHANNEL__TXDLY_LCFG_SZ 16

`define GTHE4_CHANNEL__TXDRVBIAS_N    32'h00000188
`define GTHE4_CHANNEL__TXDRVBIAS_N_SZ 4

`define GTHE4_CHANNEL__TXFIFO_ADDR_CFG    32'h00000189
`define GTHE4_CHANNEL__TXFIFO_ADDR_CFG_SZ 32

`define GTHE4_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR    32'h0000018a
`define GTHE4_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR_SZ 3

`define GTHE4_CHANNEL__TXGEARBOX_EN    32'h0000018b
`define GTHE4_CHANNEL__TXGEARBOX_EN_SZ 40

`define GTHE4_CHANNEL__TXOUT_DIV    32'h0000018c
`define GTHE4_CHANNEL__TXOUT_DIV_SZ 5

`define GTHE4_CHANNEL__TXPCSRESET_TIME    32'h0000018d
`define GTHE4_CHANNEL__TXPCSRESET_TIME_SZ 5

`define GTHE4_CHANNEL__TXPHDLY_CFG0    32'h0000018e
`define GTHE4_CHANNEL__TXPHDLY_CFG0_SZ 16

`define GTHE4_CHANNEL__TXPHDLY_CFG1    32'h0000018f
`define GTHE4_CHANNEL__TXPHDLY_CFG1_SZ 16

`define GTHE4_CHANNEL__TXPH_CFG    32'h00000190
`define GTHE4_CHANNEL__TXPH_CFG_SZ 16

`define GTHE4_CHANNEL__TXPH_CFG2    32'h00000191
`define GTHE4_CHANNEL__TXPH_CFG2_SZ 16

`define GTHE4_CHANNEL__TXPH_MONITOR_SEL    32'h00000192
`define GTHE4_CHANNEL__TXPH_MONITOR_SEL_SZ 5

`define GTHE4_CHANNEL__TXPI_CFG    32'h00000193
`define GTHE4_CHANNEL__TXPI_CFG_SZ 16

`define GTHE4_CHANNEL__TXPI_CFG0    32'h00000194
`define GTHE4_CHANNEL__TXPI_CFG0_SZ 2

`define GTHE4_CHANNEL__TXPI_CFG1    32'h00000195
`define GTHE4_CHANNEL__TXPI_CFG1_SZ 2

`define GTHE4_CHANNEL__TXPI_CFG2    32'h00000196
`define GTHE4_CHANNEL__TXPI_CFG2_SZ 2

`define GTHE4_CHANNEL__TXPI_CFG3    32'h00000197
`define GTHE4_CHANNEL__TXPI_CFG3_SZ 1

`define GTHE4_CHANNEL__TXPI_CFG4    32'h00000198
`define GTHE4_CHANNEL__TXPI_CFG4_SZ 1

`define GTHE4_CHANNEL__TXPI_CFG5    32'h00000199
`define GTHE4_CHANNEL__TXPI_CFG5_SZ 3

`define GTHE4_CHANNEL__TXPI_GRAY_SEL    32'h0000019a
`define GTHE4_CHANNEL__TXPI_GRAY_SEL_SZ 1

`define GTHE4_CHANNEL__TXPI_INVSTROBE_SEL    32'h0000019b
`define GTHE4_CHANNEL__TXPI_INVSTROBE_SEL_SZ 1

`define GTHE4_CHANNEL__TXPI_LPM    32'h0000019c
`define GTHE4_CHANNEL__TXPI_LPM_SZ 1

`define GTHE4_CHANNEL__TXPI_PPM    32'h0000019d
`define GTHE4_CHANNEL__TXPI_PPM_SZ 1

`define GTHE4_CHANNEL__TXPI_PPMCLK_SEL    32'h0000019e
`define GTHE4_CHANNEL__TXPI_PPMCLK_SEL_SZ 72

`define GTHE4_CHANNEL__TXPI_PPM_CFG    32'h0000019f
`define GTHE4_CHANNEL__TXPI_PPM_CFG_SZ 8

`define GTHE4_CHANNEL__TXPI_SYNFREQ_PPM    32'h000001a0
`define GTHE4_CHANNEL__TXPI_SYNFREQ_PPM_SZ 3

`define GTHE4_CHANNEL__TXPI_VREFSEL    32'h000001a1
`define GTHE4_CHANNEL__TXPI_VREFSEL_SZ 1

`define GTHE4_CHANNEL__TXPMARESET_TIME    32'h000001a2
`define GTHE4_CHANNEL__TXPMARESET_TIME_SZ 5

`define GTHE4_CHANNEL__TXREFCLKDIV2_SEL    32'h000001a3
`define GTHE4_CHANNEL__TXREFCLKDIV2_SEL_SZ 1

`define GTHE4_CHANNEL__TXSYNC_MULTILANE    32'h000001a4
`define GTHE4_CHANNEL__TXSYNC_MULTILANE_SZ 1

`define GTHE4_CHANNEL__TXSYNC_OVRD    32'h000001a5
`define GTHE4_CHANNEL__TXSYNC_OVRD_SZ 1

`define GTHE4_CHANNEL__TXSYNC_SKIP_DA    32'h000001a6
`define GTHE4_CHANNEL__TXSYNC_SKIP_DA_SZ 1

`define GTHE4_CHANNEL__TX_CLK25_DIV    32'h000001a7
`define GTHE4_CHANNEL__TX_CLK25_DIV_SZ 6

`define GTHE4_CHANNEL__TX_CLKMUX_EN    32'h000001a8
`define GTHE4_CHANNEL__TX_CLKMUX_EN_SZ 1

`define GTHE4_CHANNEL__TX_DATA_WIDTH    32'h000001a9
`define GTHE4_CHANNEL__TX_DATA_WIDTH_SZ 8

`define GTHE4_CHANNEL__TX_DCC_LOOP_RST_CFG    32'h000001aa
`define GTHE4_CHANNEL__TX_DCC_LOOP_RST_CFG_SZ 16

`define GTHE4_CHANNEL__TX_DEEMPH0    32'h000001ab
`define GTHE4_CHANNEL__TX_DEEMPH0_SZ 6

`define GTHE4_CHANNEL__TX_DEEMPH1    32'h000001ac
`define GTHE4_CHANNEL__TX_DEEMPH1_SZ 6

`define GTHE4_CHANNEL__TX_DEEMPH2    32'h000001ad
`define GTHE4_CHANNEL__TX_DEEMPH2_SZ 6

`define GTHE4_CHANNEL__TX_DEEMPH3    32'h000001ae
`define GTHE4_CHANNEL__TX_DEEMPH3_SZ 6

`define GTHE4_CHANNEL__TX_DIVRESET_TIME    32'h000001af
`define GTHE4_CHANNEL__TX_DIVRESET_TIME_SZ 5

`define GTHE4_CHANNEL__TX_DRIVE_MODE    32'h000001b0
`define GTHE4_CHANNEL__TX_DRIVE_MODE_SZ 64

`define GTHE4_CHANNEL__TX_DRVMUX_CTRL    32'h000001b1
`define GTHE4_CHANNEL__TX_DRVMUX_CTRL_SZ 2

`define GTHE4_CHANNEL__TX_EIDLE_ASSERT_DELAY    32'h000001b2
`define GTHE4_CHANNEL__TX_EIDLE_ASSERT_DELAY_SZ 3

`define GTHE4_CHANNEL__TX_EIDLE_DEASSERT_DELAY    32'h000001b3
`define GTHE4_CHANNEL__TX_EIDLE_DEASSERT_DELAY_SZ 3

`define GTHE4_CHANNEL__TX_FABINT_USRCLK_FLOP    32'h000001b4
`define GTHE4_CHANNEL__TX_FABINT_USRCLK_FLOP_SZ 1

`define GTHE4_CHANNEL__TX_FIFO_BYP_EN    32'h000001b5
`define GTHE4_CHANNEL__TX_FIFO_BYP_EN_SZ 1

`define GTHE4_CHANNEL__TX_IDLE_DATA_ZERO    32'h000001b6
`define GTHE4_CHANNEL__TX_IDLE_DATA_ZERO_SZ 1

`define GTHE4_CHANNEL__TX_INT_DATAWIDTH    32'h000001b7
`define GTHE4_CHANNEL__TX_INT_DATAWIDTH_SZ 2

`define GTHE4_CHANNEL__TX_LOOPBACK_DRIVE_HIZ    32'h000001b8
`define GTHE4_CHANNEL__TX_LOOPBACK_DRIVE_HIZ_SZ 40

`define GTHE4_CHANNEL__TX_MAINCURSOR_SEL    32'h000001b9
`define GTHE4_CHANNEL__TX_MAINCURSOR_SEL_SZ 1

`define GTHE4_CHANNEL__TX_MARGIN_FULL_0    32'h000001ba
`define GTHE4_CHANNEL__TX_MARGIN_FULL_0_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_FULL_1    32'h000001bb
`define GTHE4_CHANNEL__TX_MARGIN_FULL_1_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_FULL_2    32'h000001bc
`define GTHE4_CHANNEL__TX_MARGIN_FULL_2_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_FULL_3    32'h000001bd
`define GTHE4_CHANNEL__TX_MARGIN_FULL_3_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_FULL_4    32'h000001be
`define GTHE4_CHANNEL__TX_MARGIN_FULL_4_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_LOW_0    32'h000001bf
`define GTHE4_CHANNEL__TX_MARGIN_LOW_0_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_LOW_1    32'h000001c0
`define GTHE4_CHANNEL__TX_MARGIN_LOW_1_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_LOW_2    32'h000001c1
`define GTHE4_CHANNEL__TX_MARGIN_LOW_2_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_LOW_3    32'h000001c2
`define GTHE4_CHANNEL__TX_MARGIN_LOW_3_SZ 7

`define GTHE4_CHANNEL__TX_MARGIN_LOW_4    32'h000001c3
`define GTHE4_CHANNEL__TX_MARGIN_LOW_4_SZ 7

`define GTHE4_CHANNEL__TX_PHICAL_CFG0    32'h000001c4
`define GTHE4_CHANNEL__TX_PHICAL_CFG0_SZ 16

`define GTHE4_CHANNEL__TX_PHICAL_CFG1    32'h000001c5
`define GTHE4_CHANNEL__TX_PHICAL_CFG1_SZ 16

`define GTHE4_CHANNEL__TX_PHICAL_CFG2    32'h000001c6
`define GTHE4_CHANNEL__TX_PHICAL_CFG2_SZ 16

`define GTHE4_CHANNEL__TX_PI_BIASSET    32'h000001c7
`define GTHE4_CHANNEL__TX_PI_BIASSET_SZ 2

`define GTHE4_CHANNEL__TX_PI_IBIAS_MID    32'h000001c8
`define GTHE4_CHANNEL__TX_PI_IBIAS_MID_SZ 2

`define GTHE4_CHANNEL__TX_PMADATA_OPT    32'h000001c9
`define GTHE4_CHANNEL__TX_PMADATA_OPT_SZ 1

`define GTHE4_CHANNEL__TX_PMA_POWER_SAVE    32'h000001ca
`define GTHE4_CHANNEL__TX_PMA_POWER_SAVE_SZ 1

`define GTHE4_CHANNEL__TX_PMA_RSV0    32'h000001cb
`define GTHE4_CHANNEL__TX_PMA_RSV0_SZ 16

`define GTHE4_CHANNEL__TX_PREDRV_CTRL    32'h000001cc
`define GTHE4_CHANNEL__TX_PREDRV_CTRL_SZ 2

`define GTHE4_CHANNEL__TX_PROGCLK_SEL    32'h000001cd
`define GTHE4_CHANNEL__TX_PROGCLK_SEL_SZ 48

`define GTHE4_CHANNEL__TX_PROGDIV_CFG    32'h000001ce
`define GTHE4_CHANNEL__TX_PROGDIV_CFG_SZ 64

`define GTHE4_CHANNEL__TX_PROGDIV_RATE    32'h000001cf
`define GTHE4_CHANNEL__TX_PROGDIV_RATE_SZ 16

`define GTHE4_CHANNEL__TX_QPI_STATUS_EN    32'h000001d0
`define GTHE4_CHANNEL__TX_QPI_STATUS_EN_SZ 1

`define GTHE4_CHANNEL__TX_RXDETECT_CFG    32'h000001d1
`define GTHE4_CHANNEL__TX_RXDETECT_CFG_SZ 14

`define GTHE4_CHANNEL__TX_RXDETECT_REF    32'h000001d2
`define GTHE4_CHANNEL__TX_RXDETECT_REF_SZ 3

`define GTHE4_CHANNEL__TX_SAMPLE_PERIOD    32'h000001d3
`define GTHE4_CHANNEL__TX_SAMPLE_PERIOD_SZ 3

`define GTHE4_CHANNEL__TX_SARC_LPBK_ENB    32'h000001d4
`define GTHE4_CHANNEL__TX_SARC_LPBK_ENB_SZ 1

`define GTHE4_CHANNEL__TX_SW_MEAS    32'h000001d5
`define GTHE4_CHANNEL__TX_SW_MEAS_SZ 2

`define GTHE4_CHANNEL__TX_VREG_CTRL    32'h000001d6
`define GTHE4_CHANNEL__TX_VREG_CTRL_SZ 3

`define GTHE4_CHANNEL__TX_VREG_PDB    32'h000001d7
`define GTHE4_CHANNEL__TX_VREG_PDB_SZ 1

`define GTHE4_CHANNEL__TX_VREG_VREFSEL    32'h000001d8
`define GTHE4_CHANNEL__TX_VREG_VREFSEL_SZ 2

`define GTHE4_CHANNEL__TX_XCLK_SEL    32'h000001d9
`define GTHE4_CHANNEL__TX_XCLK_SEL_SZ 40

`define GTHE4_CHANNEL__USB_BOTH_BURST_IDLE    32'h000001da
`define GTHE4_CHANNEL__USB_BOTH_BURST_IDLE_SZ 1

`define GTHE4_CHANNEL__USB_BURSTMAX_U3WAKE    32'h000001db
`define GTHE4_CHANNEL__USB_BURSTMAX_U3WAKE_SZ 7

`define GTHE4_CHANNEL__USB_BURSTMIN_U3WAKE    32'h000001dc
`define GTHE4_CHANNEL__USB_BURSTMIN_U3WAKE_SZ 7

`define GTHE4_CHANNEL__USB_CLK_COR_EQ_EN    32'h000001dd
`define GTHE4_CHANNEL__USB_CLK_COR_EQ_EN_SZ 1

`define GTHE4_CHANNEL__USB_EXT_CNTL    32'h000001de
`define GTHE4_CHANNEL__USB_EXT_CNTL_SZ 1

`define GTHE4_CHANNEL__USB_IDLEMAX_POLLING    32'h000001df
`define GTHE4_CHANNEL__USB_IDLEMAX_POLLING_SZ 10

`define GTHE4_CHANNEL__USB_IDLEMIN_POLLING    32'h000001e0
`define GTHE4_CHANNEL__USB_IDLEMIN_POLLING_SZ 10

`define GTHE4_CHANNEL__USB_LFPSPING_BURST    32'h000001e1
`define GTHE4_CHANNEL__USB_LFPSPING_BURST_SZ 9

`define GTHE4_CHANNEL__USB_LFPSPOLLING_BURST    32'h000001e2
`define GTHE4_CHANNEL__USB_LFPSPOLLING_BURST_SZ 9

`define GTHE4_CHANNEL__USB_LFPSPOLLING_IDLE_MS    32'h000001e3
`define GTHE4_CHANNEL__USB_LFPSPOLLING_IDLE_MS_SZ 9

`define GTHE4_CHANNEL__USB_LFPSU1EXIT_BURST    32'h000001e4
`define GTHE4_CHANNEL__USB_LFPSU1EXIT_BURST_SZ 9

`define GTHE4_CHANNEL__USB_LFPSU2LPEXIT_BURST_MS    32'h000001e5
`define GTHE4_CHANNEL__USB_LFPSU2LPEXIT_BURST_MS_SZ 9

`define GTHE4_CHANNEL__USB_LFPSU3WAKE_BURST_MS    32'h000001e6
`define GTHE4_CHANNEL__USB_LFPSU3WAKE_BURST_MS_SZ 9

`define GTHE4_CHANNEL__USB_LFPS_TPERIOD    32'h000001e7
`define GTHE4_CHANNEL__USB_LFPS_TPERIOD_SZ 4

`define GTHE4_CHANNEL__USB_LFPS_TPERIOD_ACCURATE    32'h000001e8
`define GTHE4_CHANNEL__USB_LFPS_TPERIOD_ACCURATE_SZ 1

`define GTHE4_CHANNEL__USB_MODE    32'h000001e9
`define GTHE4_CHANNEL__USB_MODE_SZ 1

`define GTHE4_CHANNEL__USB_PCIE_ERR_REP_DIS    32'h000001ea
`define GTHE4_CHANNEL__USB_PCIE_ERR_REP_DIS_SZ 1

`define GTHE4_CHANNEL__USB_PING_SATA_MAX_INIT    32'h000001eb
`define GTHE4_CHANNEL__USB_PING_SATA_MAX_INIT_SZ 6

`define GTHE4_CHANNEL__USB_PING_SATA_MIN_INIT    32'h000001ec
`define GTHE4_CHANNEL__USB_PING_SATA_MIN_INIT_SZ 6

`define GTHE4_CHANNEL__USB_POLL_SATA_MAX_BURST    32'h000001ed
`define GTHE4_CHANNEL__USB_POLL_SATA_MAX_BURST_SZ 6

`define GTHE4_CHANNEL__USB_POLL_SATA_MIN_BURST    32'h000001ee
`define GTHE4_CHANNEL__USB_POLL_SATA_MIN_BURST_SZ 6

`define GTHE4_CHANNEL__USB_RAW_ELEC    32'h000001ef
`define GTHE4_CHANNEL__USB_RAW_ELEC_SZ 1

`define GTHE4_CHANNEL__USB_RXIDLE_P0_CTRL    32'h000001f0
`define GTHE4_CHANNEL__USB_RXIDLE_P0_CTRL_SZ 1

`define GTHE4_CHANNEL__USB_TXIDLE_TUNE_ENABLE    32'h000001f1
`define GTHE4_CHANNEL__USB_TXIDLE_TUNE_ENABLE_SZ 1

`define GTHE4_CHANNEL__USB_U1_SATA_MAX_WAKE    32'h000001f2
`define GTHE4_CHANNEL__USB_U1_SATA_MAX_WAKE_SZ 6

`define GTHE4_CHANNEL__USB_U1_SATA_MIN_WAKE    32'h000001f3
`define GTHE4_CHANNEL__USB_U1_SATA_MIN_WAKE_SZ 6

`define GTHE4_CHANNEL__USB_U2_SAS_MAX_COM    32'h000001f4
`define GTHE4_CHANNEL__USB_U2_SAS_MAX_COM_SZ 7

`define GTHE4_CHANNEL__USB_U2_SAS_MIN_COM    32'h000001f5
`define GTHE4_CHANNEL__USB_U2_SAS_MIN_COM_SZ 6

`define GTHE4_CHANNEL__USE_PCS_CLK_PHASE_SEL    32'h000001f6
`define GTHE4_CHANNEL__USE_PCS_CLK_PHASE_SEL_SZ 1

`define GTHE4_CHANNEL__Y_ALL_MODE    32'h000001f7
`define GTHE4_CHANNEL__Y_ALL_MODE_SZ 1

`endif  // B_GTHE4_CHANNEL_DEFINES_VH