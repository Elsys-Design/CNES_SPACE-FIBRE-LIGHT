// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_X5PHIO_CMUIF_DEFINES_VH
`else
`define B_X5PHIO_CMUIF_DEFINES_VH

// Look-up table parameters
//

`define X5PHIO_CMUIF_ADDR_N  4
`define X5PHIO_CMUIF_ADDR_SZ 32
`define X5PHIO_CMUIF_DATA_SZ 40

// Attribute addresses
//

`define X5PHIO_CMUIF__APBCLK_FREQ    32'h00000000
`define X5PHIO_CMUIF__APBCLK_FREQ_SZ 9

`define X5PHIO_CMUIF__DMC_APB_SEL_CMU    32'h00000001
`define X5PHIO_CMUIF__DMC_APB_SEL_CMU_SZ 40

`define X5PHIO_CMUIF__RIUCLK_DBLR_BYPASS    32'h00000002
`define X5PHIO_CMUIF__RIUCLK_DBLR_BYPASS_SZ 40

`define X5PHIO_CMUIF__RIU_CLK_DBL_CMU    32'h00000003
`define X5PHIO_CMUIF__RIU_CLK_DBL_CMU_SZ 3

`endif  // B_X5PHIO_CMUIF_DEFINES_VH