// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DDRMC5_DEFINES_VH
`else
`define B_DDRMC5_DEFINES_VH

// Look-up table parameters
//

`define DDRMC5_ADDR_N  626
`define DDRMC5_ADDR_SZ 32
`define DDRMC5_DATA_SZ 32

// Attribute addresses
//

`define DDRMC5__A2A_CNTRL_MAP_0    32'h00000000
`define DDRMC5__A2A_CNTRL_MAP_0_SZ 30

`define DDRMC5__A2A_CNTRL_MAP_1    32'h00000001
`define DDRMC5__A2A_CNTRL_MAP_1_SZ 30

`define DDRMC5__A2A_CNTRL_MAP_2    32'h00000002
`define DDRMC5__A2A_CNTRL_MAP_2_SZ 12

`define DDRMC5__A2A_DIFF_C_PIN_MAP_0    32'h00000003
`define DDRMC5__A2A_DIFF_C_PIN_MAP_0_SZ 30

`define DDRMC5__A2A_DIFF_C_PIN_MAP_1    32'h00000004
`define DDRMC5__A2A_DIFF_C_PIN_MAP_1_SZ 30

`define DDRMC5__A2A_DIFF_C_PIN_MAP_2    32'h00000005
`define DDRMC5__A2A_DIFF_C_PIN_MAP_2_SZ 12

`define DDRMC5__A2A_DIFF_T_PIN_MAP_0    32'h00000006
`define DDRMC5__A2A_DIFF_T_PIN_MAP_0_SZ 30

`define DDRMC5__A2A_DIFF_T_PIN_MAP_1    32'h00000007
`define DDRMC5__A2A_DIFF_T_PIN_MAP_1_SZ 30

`define DDRMC5__A2A_DIFF_T_PIN_MAP_2    32'h00000008
`define DDRMC5__A2A_DIFF_T_PIN_MAP_2_SZ 12

`define DDRMC5__A2A_DUAL_CHAN    32'h00000009
`define DDRMC5__A2A_DUAL_CHAN_SZ 1

`define DDRMC5__A2A_PIN_MAP_0    32'h0000000a
`define DDRMC5__A2A_PIN_MAP_0_SZ 28

`define DDRMC5__A2A_PIN_MAP_1    32'h0000000b
`define DDRMC5__A2A_PIN_MAP_1_SZ 28

`define DDRMC5__A2A_PIN_MAP_10    32'h0000000c
`define DDRMC5__A2A_PIN_MAP_10_SZ 28

`define DDRMC5__A2A_PIN_MAP_11    32'h0000000d
`define DDRMC5__A2A_PIN_MAP_11_SZ 28

`define DDRMC5__A2A_PIN_MAP_12    32'h0000000e
`define DDRMC5__A2A_PIN_MAP_12_SZ 28

`define DDRMC5__A2A_PIN_MAP_13    32'h0000000f
`define DDRMC5__A2A_PIN_MAP_13_SZ 28

`define DDRMC5__A2A_PIN_MAP_14    32'h00000010
`define DDRMC5__A2A_PIN_MAP_14_SZ 28

`define DDRMC5__A2A_PIN_MAP_15    32'h00000011
`define DDRMC5__A2A_PIN_MAP_15_SZ 28

`define DDRMC5__A2A_PIN_MAP_16    32'h00000012
`define DDRMC5__A2A_PIN_MAP_16_SZ 28

`define DDRMC5__A2A_PIN_MAP_17    32'h00000013
`define DDRMC5__A2A_PIN_MAP_17_SZ 28

`define DDRMC5__A2A_PIN_MAP_2    32'h00000014
`define DDRMC5__A2A_PIN_MAP_2_SZ 28

`define DDRMC5__A2A_PIN_MAP_3    32'h00000015
`define DDRMC5__A2A_PIN_MAP_3_SZ 28

`define DDRMC5__A2A_PIN_MAP_4    32'h00000016
`define DDRMC5__A2A_PIN_MAP_4_SZ 28

`define DDRMC5__A2A_PIN_MAP_5    32'h00000017
`define DDRMC5__A2A_PIN_MAP_5_SZ 28

`define DDRMC5__A2A_PIN_MAP_6    32'h00000018
`define DDRMC5__A2A_PIN_MAP_6_SZ 28

`define DDRMC5__A2A_PIN_MAP_7    32'h00000019
`define DDRMC5__A2A_PIN_MAP_7_SZ 28

`define DDRMC5__A2A_PIN_MAP_8    32'h0000001a
`define DDRMC5__A2A_PIN_MAP_8_SZ 28

`define DDRMC5__A2A_PIN_MAP_9    32'h0000001b
`define DDRMC5__A2A_PIN_MAP_9_SZ 28

`define DDRMC5__A2A_RD_MAP    32'h0000001c
`define DDRMC5__A2A_RD_MAP_SZ 14

`define DDRMC5__A2A_RD_MAP_DBI_CH0_0    32'h0000001d
`define DDRMC5__A2A_RD_MAP_DBI_CH0_0_SZ 28

`define DDRMC5__A2A_RD_MAP_DBI_CH0_1    32'h0000001e
`define DDRMC5__A2A_RD_MAP_DBI_CH0_1_SZ 7

`define DDRMC5__A2A_RD_MAP_DBI_CH1_0    32'h0000001f
`define DDRMC5__A2A_RD_MAP_DBI_CH1_0_SZ 28

`define DDRMC5__A2A_RD_MAP_DBI_CH1_1    32'h00000020
`define DDRMC5__A2A_RD_MAP_DBI_CH1_1_SZ 7

`define DDRMC5__A2A_RD_MAP_DQ_0    32'h00000021
`define DDRMC5__A2A_RD_MAP_DQ_0_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_1    32'h00000022
`define DDRMC5__A2A_RD_MAP_DQ_1_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_2    32'h00000023
`define DDRMC5__A2A_RD_MAP_DQ_2_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_3    32'h00000024
`define DDRMC5__A2A_RD_MAP_DQ_3_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_4    32'h00000025
`define DDRMC5__A2A_RD_MAP_DQ_4_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_5    32'h00000026
`define DDRMC5__A2A_RD_MAP_DQ_5_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_6    32'h00000027
`define DDRMC5__A2A_RD_MAP_DQ_6_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_7    32'h00000028
`define DDRMC5__A2A_RD_MAP_DQ_7_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_8    32'h00000029
`define DDRMC5__A2A_RD_MAP_DQ_8_SZ 28

`define DDRMC5__A2A_RD_MAP_DQ_9    32'h0000002a
`define DDRMC5__A2A_RD_MAP_DQ_9_SZ 28

`define DDRMC5__ARBITER_CONFIG    32'h0000002b
`define DDRMC5__ARBITER_CONFIG_SZ 1

`define DDRMC5__CAL_CS_CH    32'h0000002c
`define DDRMC5__CAL_CS_CH_SZ 3

`define DDRMC5__CAL_MODE    32'h0000002d
`define DDRMC5__CAL_MODE_SZ 1

`define DDRMC5__CK_PATTERN    32'h0000002e
`define DDRMC5__CK_PATTERN_SZ 17

`define DDRMC5__CLK_GATE    32'h0000002f
`define DDRMC5__CLK_GATE_SZ 22

`define DDRMC5__CPLX_BURST_ARRAY0    32'h00000030
`define DDRMC5__CPLX_BURST_ARRAY0_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY1    32'h00000031
`define DDRMC5__CPLX_BURST_ARRAY1_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY10    32'h00000032
`define DDRMC5__CPLX_BURST_ARRAY10_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY11    32'h00000033
`define DDRMC5__CPLX_BURST_ARRAY11_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY12    32'h00000034
`define DDRMC5__CPLX_BURST_ARRAY12_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY13    32'h00000035
`define DDRMC5__CPLX_BURST_ARRAY13_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY14    32'h00000036
`define DDRMC5__CPLX_BURST_ARRAY14_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY15    32'h00000037
`define DDRMC5__CPLX_BURST_ARRAY15_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY16    32'h00000038
`define DDRMC5__CPLX_BURST_ARRAY16_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY17    32'h00000039
`define DDRMC5__CPLX_BURST_ARRAY17_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY18    32'h0000003a
`define DDRMC5__CPLX_BURST_ARRAY18_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY19    32'h0000003b
`define DDRMC5__CPLX_BURST_ARRAY19_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY2    32'h0000003c
`define DDRMC5__CPLX_BURST_ARRAY2_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY20    32'h0000003d
`define DDRMC5__CPLX_BURST_ARRAY20_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY21    32'h0000003e
`define DDRMC5__CPLX_BURST_ARRAY21_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY22    32'h0000003f
`define DDRMC5__CPLX_BURST_ARRAY22_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY3    32'h00000040
`define DDRMC5__CPLX_BURST_ARRAY3_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY4    32'h00000041
`define DDRMC5__CPLX_BURST_ARRAY4_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY5    32'h00000042
`define DDRMC5__CPLX_BURST_ARRAY5_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY6    32'h00000043
`define DDRMC5__CPLX_BURST_ARRAY6_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY7    32'h00000044
`define DDRMC5__CPLX_BURST_ARRAY7_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY8    32'h00000045
`define DDRMC5__CPLX_BURST_ARRAY8_SZ 5

`define DDRMC5__CPLX_BURST_ARRAY9    32'h00000046
`define DDRMC5__CPLX_BURST_ARRAY9_SZ 5

`define DDRMC5__CPLX_CONFIG2    32'h00000047
`define DDRMC5__CPLX_CONFIG2_SZ 25

`define DDRMC5__CPLX_PATTERN0    32'h00000048
`define DDRMC5__CPLX_PATTERN0_SZ 16

`define DDRMC5__CPLX_PATTERN1    32'h00000049
`define DDRMC5__CPLX_PATTERN1_SZ 16

`define DDRMC5__CPLX_PATTERN10    32'h0000004a
`define DDRMC5__CPLX_PATTERN10_SZ 16

`define DDRMC5__CPLX_PATTERN100    32'h0000004b
`define DDRMC5__CPLX_PATTERN100_SZ 16

`define DDRMC5__CPLX_PATTERN101    32'h0000004c
`define DDRMC5__CPLX_PATTERN101_SZ 16

`define DDRMC5__CPLX_PATTERN102    32'h0000004d
`define DDRMC5__CPLX_PATTERN102_SZ 16

`define DDRMC5__CPLX_PATTERN103    32'h0000004e
`define DDRMC5__CPLX_PATTERN103_SZ 16

`define DDRMC5__CPLX_PATTERN104    32'h0000004f
`define DDRMC5__CPLX_PATTERN104_SZ 16

`define DDRMC5__CPLX_PATTERN105    32'h00000050
`define DDRMC5__CPLX_PATTERN105_SZ 16

`define DDRMC5__CPLX_PATTERN106    32'h00000051
`define DDRMC5__CPLX_PATTERN106_SZ 16

`define DDRMC5__CPLX_PATTERN107    32'h00000052
`define DDRMC5__CPLX_PATTERN107_SZ 16

`define DDRMC5__CPLX_PATTERN108    32'h00000053
`define DDRMC5__CPLX_PATTERN108_SZ 16

`define DDRMC5__CPLX_PATTERN109    32'h00000054
`define DDRMC5__CPLX_PATTERN109_SZ 16

`define DDRMC5__CPLX_PATTERN11    32'h00000055
`define DDRMC5__CPLX_PATTERN11_SZ 16

`define DDRMC5__CPLX_PATTERN110    32'h00000056
`define DDRMC5__CPLX_PATTERN110_SZ 16

`define DDRMC5__CPLX_PATTERN111    32'h00000057
`define DDRMC5__CPLX_PATTERN111_SZ 16

`define DDRMC5__CPLX_PATTERN112    32'h00000058
`define DDRMC5__CPLX_PATTERN112_SZ 16

`define DDRMC5__CPLX_PATTERN113    32'h00000059
`define DDRMC5__CPLX_PATTERN113_SZ 16

`define DDRMC5__CPLX_PATTERN114    32'h0000005a
`define DDRMC5__CPLX_PATTERN114_SZ 16

`define DDRMC5__CPLX_PATTERN115    32'h0000005b
`define DDRMC5__CPLX_PATTERN115_SZ 16

`define DDRMC5__CPLX_PATTERN116    32'h0000005c
`define DDRMC5__CPLX_PATTERN116_SZ 16

`define DDRMC5__CPLX_PATTERN117    32'h0000005d
`define DDRMC5__CPLX_PATTERN117_SZ 16

`define DDRMC5__CPLX_PATTERN118    32'h0000005e
`define DDRMC5__CPLX_PATTERN118_SZ 16

`define DDRMC5__CPLX_PATTERN119    32'h0000005f
`define DDRMC5__CPLX_PATTERN119_SZ 16

`define DDRMC5__CPLX_PATTERN12    32'h00000060
`define DDRMC5__CPLX_PATTERN12_SZ 16

`define DDRMC5__CPLX_PATTERN120    32'h00000061
`define DDRMC5__CPLX_PATTERN120_SZ 16

`define DDRMC5__CPLX_PATTERN121    32'h00000062
`define DDRMC5__CPLX_PATTERN121_SZ 16

`define DDRMC5__CPLX_PATTERN122    32'h00000063
`define DDRMC5__CPLX_PATTERN122_SZ 16

`define DDRMC5__CPLX_PATTERN123    32'h00000064
`define DDRMC5__CPLX_PATTERN123_SZ 16

`define DDRMC5__CPLX_PATTERN124    32'h00000065
`define DDRMC5__CPLX_PATTERN124_SZ 16

`define DDRMC5__CPLX_PATTERN125    32'h00000066
`define DDRMC5__CPLX_PATTERN125_SZ 16

`define DDRMC5__CPLX_PATTERN126    32'h00000067
`define DDRMC5__CPLX_PATTERN126_SZ 16

`define DDRMC5__CPLX_PATTERN127    32'h00000068
`define DDRMC5__CPLX_PATTERN127_SZ 16

`define DDRMC5__CPLX_PATTERN128    32'h00000069
`define DDRMC5__CPLX_PATTERN128_SZ 16

`define DDRMC5__CPLX_PATTERN129    32'h0000006a
`define DDRMC5__CPLX_PATTERN129_SZ 16

`define DDRMC5__CPLX_PATTERN13    32'h0000006b
`define DDRMC5__CPLX_PATTERN13_SZ 16

`define DDRMC5__CPLX_PATTERN130    32'h0000006c
`define DDRMC5__CPLX_PATTERN130_SZ 16

`define DDRMC5__CPLX_PATTERN131    32'h0000006d
`define DDRMC5__CPLX_PATTERN131_SZ 16

`define DDRMC5__CPLX_PATTERN132    32'h0000006e
`define DDRMC5__CPLX_PATTERN132_SZ 16

`define DDRMC5__CPLX_PATTERN133    32'h0000006f
`define DDRMC5__CPLX_PATTERN133_SZ 16

`define DDRMC5__CPLX_PATTERN134    32'h00000070
`define DDRMC5__CPLX_PATTERN134_SZ 16

`define DDRMC5__CPLX_PATTERN135    32'h00000071
`define DDRMC5__CPLX_PATTERN135_SZ 16

`define DDRMC5__CPLX_PATTERN136    32'h00000072
`define DDRMC5__CPLX_PATTERN136_SZ 16

`define DDRMC5__CPLX_PATTERN137    32'h00000073
`define DDRMC5__CPLX_PATTERN137_SZ 16

`define DDRMC5__CPLX_PATTERN138    32'h00000074
`define DDRMC5__CPLX_PATTERN138_SZ 16

`define DDRMC5__CPLX_PATTERN139    32'h00000075
`define DDRMC5__CPLX_PATTERN139_SZ 16

`define DDRMC5__CPLX_PATTERN14    32'h00000076
`define DDRMC5__CPLX_PATTERN14_SZ 16

`define DDRMC5__CPLX_PATTERN140    32'h00000077
`define DDRMC5__CPLX_PATTERN140_SZ 16

`define DDRMC5__CPLX_PATTERN141    32'h00000078
`define DDRMC5__CPLX_PATTERN141_SZ 16

`define DDRMC5__CPLX_PATTERN142    32'h00000079
`define DDRMC5__CPLX_PATTERN142_SZ 16

`define DDRMC5__CPLX_PATTERN143    32'h0000007a
`define DDRMC5__CPLX_PATTERN143_SZ 16

`define DDRMC5__CPLX_PATTERN144    32'h0000007b
`define DDRMC5__CPLX_PATTERN144_SZ 16

`define DDRMC5__CPLX_PATTERN145    32'h0000007c
`define DDRMC5__CPLX_PATTERN145_SZ 16

`define DDRMC5__CPLX_PATTERN146    32'h0000007d
`define DDRMC5__CPLX_PATTERN146_SZ 16

`define DDRMC5__CPLX_PATTERN147    32'h0000007e
`define DDRMC5__CPLX_PATTERN147_SZ 16

`define DDRMC5__CPLX_PATTERN148    32'h0000007f
`define DDRMC5__CPLX_PATTERN148_SZ 16

`define DDRMC5__CPLX_PATTERN149    32'h00000080
`define DDRMC5__CPLX_PATTERN149_SZ 16

`define DDRMC5__CPLX_PATTERN15    32'h00000081
`define DDRMC5__CPLX_PATTERN15_SZ 16

`define DDRMC5__CPLX_PATTERN150    32'h00000082
`define DDRMC5__CPLX_PATTERN150_SZ 16

`define DDRMC5__CPLX_PATTERN151    32'h00000083
`define DDRMC5__CPLX_PATTERN151_SZ 16

`define DDRMC5__CPLX_PATTERN152    32'h00000084
`define DDRMC5__CPLX_PATTERN152_SZ 16

`define DDRMC5__CPLX_PATTERN153    32'h00000085
`define DDRMC5__CPLX_PATTERN153_SZ 16

`define DDRMC5__CPLX_PATTERN154    32'h00000086
`define DDRMC5__CPLX_PATTERN154_SZ 16

`define DDRMC5__CPLX_PATTERN155    32'h00000087
`define DDRMC5__CPLX_PATTERN155_SZ 16

`define DDRMC5__CPLX_PATTERN156    32'h00000088
`define DDRMC5__CPLX_PATTERN156_SZ 16

`define DDRMC5__CPLX_PATTERN16    32'h00000089
`define DDRMC5__CPLX_PATTERN16_SZ 16

`define DDRMC5__CPLX_PATTERN17    32'h0000008a
`define DDRMC5__CPLX_PATTERN17_SZ 16

`define DDRMC5__CPLX_PATTERN18    32'h0000008b
`define DDRMC5__CPLX_PATTERN18_SZ 16

`define DDRMC5__CPLX_PATTERN19    32'h0000008c
`define DDRMC5__CPLX_PATTERN19_SZ 16

`define DDRMC5__CPLX_PATTERN2    32'h0000008d
`define DDRMC5__CPLX_PATTERN2_SZ 16

`define DDRMC5__CPLX_PATTERN20    32'h0000008e
`define DDRMC5__CPLX_PATTERN20_SZ 16

`define DDRMC5__CPLX_PATTERN21    32'h0000008f
`define DDRMC5__CPLX_PATTERN21_SZ 16

`define DDRMC5__CPLX_PATTERN22    32'h00000090
`define DDRMC5__CPLX_PATTERN22_SZ 16

`define DDRMC5__CPLX_PATTERN23    32'h00000091
`define DDRMC5__CPLX_PATTERN23_SZ 16

`define DDRMC5__CPLX_PATTERN24    32'h00000092
`define DDRMC5__CPLX_PATTERN24_SZ 16

`define DDRMC5__CPLX_PATTERN25    32'h00000093
`define DDRMC5__CPLX_PATTERN25_SZ 16

`define DDRMC5__CPLX_PATTERN26    32'h00000094
`define DDRMC5__CPLX_PATTERN26_SZ 16

`define DDRMC5__CPLX_PATTERN27    32'h00000095
`define DDRMC5__CPLX_PATTERN27_SZ 16

`define DDRMC5__CPLX_PATTERN28    32'h00000096
`define DDRMC5__CPLX_PATTERN28_SZ 16

`define DDRMC5__CPLX_PATTERN29    32'h00000097
`define DDRMC5__CPLX_PATTERN29_SZ 16

`define DDRMC5__CPLX_PATTERN3    32'h00000098
`define DDRMC5__CPLX_PATTERN3_SZ 16

`define DDRMC5__CPLX_PATTERN30    32'h00000099
`define DDRMC5__CPLX_PATTERN30_SZ 16

`define DDRMC5__CPLX_PATTERN31    32'h0000009a
`define DDRMC5__CPLX_PATTERN31_SZ 16

`define DDRMC5__CPLX_PATTERN32    32'h0000009b
`define DDRMC5__CPLX_PATTERN32_SZ 16

`define DDRMC5__CPLX_PATTERN33    32'h0000009c
`define DDRMC5__CPLX_PATTERN33_SZ 16

`define DDRMC5__CPLX_PATTERN34    32'h0000009d
`define DDRMC5__CPLX_PATTERN34_SZ 16

`define DDRMC5__CPLX_PATTERN35    32'h0000009e
`define DDRMC5__CPLX_PATTERN35_SZ 16

`define DDRMC5__CPLX_PATTERN36    32'h0000009f
`define DDRMC5__CPLX_PATTERN36_SZ 16

`define DDRMC5__CPLX_PATTERN37    32'h000000a0
`define DDRMC5__CPLX_PATTERN37_SZ 16

`define DDRMC5__CPLX_PATTERN38    32'h000000a1
`define DDRMC5__CPLX_PATTERN38_SZ 16

`define DDRMC5__CPLX_PATTERN39    32'h000000a2
`define DDRMC5__CPLX_PATTERN39_SZ 16

`define DDRMC5__CPLX_PATTERN4    32'h000000a3
`define DDRMC5__CPLX_PATTERN4_SZ 16

`define DDRMC5__CPLX_PATTERN40    32'h000000a4
`define DDRMC5__CPLX_PATTERN40_SZ 16

`define DDRMC5__CPLX_PATTERN41    32'h000000a5
`define DDRMC5__CPLX_PATTERN41_SZ 16

`define DDRMC5__CPLX_PATTERN42    32'h000000a6
`define DDRMC5__CPLX_PATTERN42_SZ 16

`define DDRMC5__CPLX_PATTERN43    32'h000000a7
`define DDRMC5__CPLX_PATTERN43_SZ 16

`define DDRMC5__CPLX_PATTERN44    32'h000000a8
`define DDRMC5__CPLX_PATTERN44_SZ 16

`define DDRMC5__CPLX_PATTERN45    32'h000000a9
`define DDRMC5__CPLX_PATTERN45_SZ 16

`define DDRMC5__CPLX_PATTERN46    32'h000000aa
`define DDRMC5__CPLX_PATTERN46_SZ 16

`define DDRMC5__CPLX_PATTERN47    32'h000000ab
`define DDRMC5__CPLX_PATTERN47_SZ 16

`define DDRMC5__CPLX_PATTERN48    32'h000000ac
`define DDRMC5__CPLX_PATTERN48_SZ 16

`define DDRMC5__CPLX_PATTERN49    32'h000000ad
`define DDRMC5__CPLX_PATTERN49_SZ 16

`define DDRMC5__CPLX_PATTERN5    32'h000000ae
`define DDRMC5__CPLX_PATTERN5_SZ 16

`define DDRMC5__CPLX_PATTERN50    32'h000000af
`define DDRMC5__CPLX_PATTERN50_SZ 16

`define DDRMC5__CPLX_PATTERN51    32'h000000b0
`define DDRMC5__CPLX_PATTERN51_SZ 16

`define DDRMC5__CPLX_PATTERN52    32'h000000b1
`define DDRMC5__CPLX_PATTERN52_SZ 16

`define DDRMC5__CPLX_PATTERN53    32'h000000b2
`define DDRMC5__CPLX_PATTERN53_SZ 16

`define DDRMC5__CPLX_PATTERN54    32'h000000b3
`define DDRMC5__CPLX_PATTERN54_SZ 16

`define DDRMC5__CPLX_PATTERN55    32'h000000b4
`define DDRMC5__CPLX_PATTERN55_SZ 16

`define DDRMC5__CPLX_PATTERN56    32'h000000b5
`define DDRMC5__CPLX_PATTERN56_SZ 16

`define DDRMC5__CPLX_PATTERN57    32'h000000b6
`define DDRMC5__CPLX_PATTERN57_SZ 16

`define DDRMC5__CPLX_PATTERN58    32'h000000b7
`define DDRMC5__CPLX_PATTERN58_SZ 16

`define DDRMC5__CPLX_PATTERN59    32'h000000b8
`define DDRMC5__CPLX_PATTERN59_SZ 16

`define DDRMC5__CPLX_PATTERN6    32'h000000b9
`define DDRMC5__CPLX_PATTERN6_SZ 16

`define DDRMC5__CPLX_PATTERN60    32'h000000ba
`define DDRMC5__CPLX_PATTERN60_SZ 16

`define DDRMC5__CPLX_PATTERN61    32'h000000bb
`define DDRMC5__CPLX_PATTERN61_SZ 16

`define DDRMC5__CPLX_PATTERN62    32'h000000bc
`define DDRMC5__CPLX_PATTERN62_SZ 16

`define DDRMC5__CPLX_PATTERN63    32'h000000bd
`define DDRMC5__CPLX_PATTERN63_SZ 16

`define DDRMC5__CPLX_PATTERN64    32'h000000be
`define DDRMC5__CPLX_PATTERN64_SZ 16

`define DDRMC5__CPLX_PATTERN65    32'h000000bf
`define DDRMC5__CPLX_PATTERN65_SZ 16

`define DDRMC5__CPLX_PATTERN66    32'h000000c0
`define DDRMC5__CPLX_PATTERN66_SZ 16

`define DDRMC5__CPLX_PATTERN67    32'h000000c1
`define DDRMC5__CPLX_PATTERN67_SZ 16

`define DDRMC5__CPLX_PATTERN68    32'h000000c2
`define DDRMC5__CPLX_PATTERN68_SZ 16

`define DDRMC5__CPLX_PATTERN69    32'h000000c3
`define DDRMC5__CPLX_PATTERN69_SZ 16

`define DDRMC5__CPLX_PATTERN7    32'h000000c4
`define DDRMC5__CPLX_PATTERN7_SZ 16

`define DDRMC5__CPLX_PATTERN70    32'h000000c5
`define DDRMC5__CPLX_PATTERN70_SZ 16

`define DDRMC5__CPLX_PATTERN71    32'h000000c6
`define DDRMC5__CPLX_PATTERN71_SZ 16

`define DDRMC5__CPLX_PATTERN72    32'h000000c7
`define DDRMC5__CPLX_PATTERN72_SZ 16

`define DDRMC5__CPLX_PATTERN73    32'h000000c8
`define DDRMC5__CPLX_PATTERN73_SZ 16

`define DDRMC5__CPLX_PATTERN74    32'h000000c9
`define DDRMC5__CPLX_PATTERN74_SZ 16

`define DDRMC5__CPLX_PATTERN75    32'h000000ca
`define DDRMC5__CPLX_PATTERN75_SZ 16

`define DDRMC5__CPLX_PATTERN76    32'h000000cb
`define DDRMC5__CPLX_PATTERN76_SZ 16

`define DDRMC5__CPLX_PATTERN77    32'h000000cc
`define DDRMC5__CPLX_PATTERN77_SZ 16

`define DDRMC5__CPLX_PATTERN78    32'h000000cd
`define DDRMC5__CPLX_PATTERN78_SZ 16

`define DDRMC5__CPLX_PATTERN79    32'h000000ce
`define DDRMC5__CPLX_PATTERN79_SZ 16

`define DDRMC5__CPLX_PATTERN8    32'h000000cf
`define DDRMC5__CPLX_PATTERN8_SZ 16

`define DDRMC5__CPLX_PATTERN80    32'h000000d0
`define DDRMC5__CPLX_PATTERN80_SZ 16

`define DDRMC5__CPLX_PATTERN81    32'h000000d1
`define DDRMC5__CPLX_PATTERN81_SZ 16

`define DDRMC5__CPLX_PATTERN82    32'h000000d2
`define DDRMC5__CPLX_PATTERN82_SZ 16

`define DDRMC5__CPLX_PATTERN83    32'h000000d3
`define DDRMC5__CPLX_PATTERN83_SZ 16

`define DDRMC5__CPLX_PATTERN84    32'h000000d4
`define DDRMC5__CPLX_PATTERN84_SZ 16

`define DDRMC5__CPLX_PATTERN85    32'h000000d5
`define DDRMC5__CPLX_PATTERN85_SZ 16

`define DDRMC5__CPLX_PATTERN86    32'h000000d6
`define DDRMC5__CPLX_PATTERN86_SZ 16

`define DDRMC5__CPLX_PATTERN87    32'h000000d7
`define DDRMC5__CPLX_PATTERN87_SZ 16

`define DDRMC5__CPLX_PATTERN88    32'h000000d8
`define DDRMC5__CPLX_PATTERN88_SZ 16

`define DDRMC5__CPLX_PATTERN89    32'h000000d9
`define DDRMC5__CPLX_PATTERN89_SZ 16

`define DDRMC5__CPLX_PATTERN9    32'h000000da
`define DDRMC5__CPLX_PATTERN9_SZ 16

`define DDRMC5__CPLX_PATTERN90    32'h000000db
`define DDRMC5__CPLX_PATTERN90_SZ 16

`define DDRMC5__CPLX_PATTERN91    32'h000000dc
`define DDRMC5__CPLX_PATTERN91_SZ 16

`define DDRMC5__CPLX_PATTERN92    32'h000000dd
`define DDRMC5__CPLX_PATTERN92_SZ 16

`define DDRMC5__CPLX_PATTERN93    32'h000000de
`define DDRMC5__CPLX_PATTERN93_SZ 16

`define DDRMC5__CPLX_PATTERN94    32'h000000df
`define DDRMC5__CPLX_PATTERN94_SZ 16

`define DDRMC5__CPLX_PATTERN95    32'h000000e0
`define DDRMC5__CPLX_PATTERN95_SZ 16

`define DDRMC5__CPLX_PATTERN96    32'h000000e1
`define DDRMC5__CPLX_PATTERN96_SZ 16

`define DDRMC5__CPLX_PATTERN97    32'h000000e2
`define DDRMC5__CPLX_PATTERN97_SZ 16

`define DDRMC5__CPLX_PATTERN98    32'h000000e3
`define DDRMC5__CPLX_PATTERN98_SZ 16

`define DDRMC5__CPLX_PATTERN99    32'h000000e4
`define DDRMC5__CPLX_PATTERN99_SZ 16

`define DDRMC5__CRYPTO_TRSS_CONFIG    32'h000000e5
`define DDRMC5__CRYPTO_TRSS_CONFIG_SZ 32

`define DDRMC5__CRYPTO_TRSS_CONFIG2    32'h000000e6
`define DDRMC5__CRYPTO_TRSS_CONFIG2_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR0    32'h000000e7
`define DDRMC5__CRYPTO_TRSS_PSTR0_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR1    32'h000000e8
`define DDRMC5__CRYPTO_TRSS_PSTR1_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR10    32'h000000e9
`define DDRMC5__CRYPTO_TRSS_PSTR10_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR11    32'h000000ea
`define DDRMC5__CRYPTO_TRSS_PSTR11_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR2    32'h000000eb
`define DDRMC5__CRYPTO_TRSS_PSTR2_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR3    32'h000000ec
`define DDRMC5__CRYPTO_TRSS_PSTR3_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR4    32'h000000ed
`define DDRMC5__CRYPTO_TRSS_PSTR4_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR5    32'h000000ee
`define DDRMC5__CRYPTO_TRSS_PSTR5_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR6    32'h000000ef
`define DDRMC5__CRYPTO_TRSS_PSTR6_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR7    32'h000000f0
`define DDRMC5__CRYPTO_TRSS_PSTR7_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR8    32'h000000f1
`define DDRMC5__CRYPTO_TRSS_PSTR8_SZ 32

`define DDRMC5__CRYPTO_TRSS_PSTR9    32'h000000f2
`define DDRMC5__CRYPTO_TRSS_PSTR9_SZ 32

`define DDRMC5__DBG_TRIGGER    32'h000000f3
`define DDRMC5__DBG_TRIGGER_SZ 3

`define DDRMC5__DDR5_READ_LFSR_CFG    32'h000000f4
`define DDRMC5__DDR5_READ_LFSR_CFG_SZ 17

`define DDRMC5__DDR5_READ_LFSR_INVERT_31_0    32'h000000f5
`define DDRMC5__DDR5_READ_LFSR_INVERT_31_0_SZ 32

`define DDRMC5__DDR5_READ_LFSR_INVERT_39_32    32'h000000f6
`define DDRMC5__DDR5_READ_LFSR_INVERT_39_32_SZ 8

`define DDRMC5__DDR5_READ_LFSR_OPT_31_0    32'h000000f7
`define DDRMC5__DDR5_READ_LFSR_OPT_31_0_SZ 32

`define DDRMC5__DDR5_READ_LFSR_OPT_39_32    32'h000000f8
`define DDRMC5__DDR5_READ_LFSR_OPT_39_32_SZ 8

`define DDRMC5__DDR5_READ_LFSR_PAT_31_0    32'h000000f9
`define DDRMC5__DDR5_READ_LFSR_PAT_31_0_SZ 32

`define DDRMC5__DDR5_READ_LFSR_PAT_39_32    32'h000000fa
`define DDRMC5__DDR5_READ_LFSR_PAT_39_32_SZ 8

`define DDRMC5__DDR5_SPARE_DYN_CFG0    32'h000000fb
`define DDRMC5__DDR5_SPARE_DYN_CFG0_SZ 32

`define DDRMC5__DDR5_SPARE_STA_CFG0    32'h000000fc
`define DDRMC5__DDR5_SPARE_STA_CFG0_SZ 32

`define DDRMC5__EXMON_CLR_EXE    32'h000000fd
`define DDRMC5__EXMON_CLR_EXE_SZ 9

`define DDRMC5__FIFO_RDEN    32'h000000fe
`define DDRMC5__FIFO_RDEN_SZ 7

`define DDRMC5__LP5_MRS_BIT_MUX_BYTE0    32'h000000ff
`define DDRMC5__LP5_MRS_BIT_MUX_BYTE0_SZ 24

`define DDRMC5__LP5_MRS_BIT_MUX_BYTE1    32'h00000100
`define DDRMC5__LP5_MRS_BIT_MUX_BYTE1_SZ 24

`define DDRMC5__LP5_MRS_BIT_MUX_BYTE2    32'h00000101
`define DDRMC5__LP5_MRS_BIT_MUX_BYTE2_SZ 24

`define DDRMC5__LP5_MRS_BIT_MUX_BYTE3    32'h00000102
`define DDRMC5__LP5_MRS_BIT_MUX_BYTE3_SZ 24

`define DDRMC5__PHY_RANK_READ_OVERRIDE    32'h00000103
`define DDRMC5__PHY_RANK_READ_OVERRIDE_SZ 18

`define DDRMC5__PHY_RANK_WRITE_OVERRIDE    32'h00000104
`define DDRMC5__PHY_RANK_WRITE_OVERRIDE_SZ 18

`define DDRMC5__PHY_RDEN0    32'h00000105
`define DDRMC5__PHY_RDEN0_SZ 8

`define DDRMC5__PHY_RDEN1    32'h00000106
`define DDRMC5__PHY_RDEN1_SZ 8

`define DDRMC5__PHY_RDEN2    32'h00000107
`define DDRMC5__PHY_RDEN2_SZ 8

`define DDRMC5__PHY_RDEN3    32'h00000108
`define DDRMC5__PHY_RDEN3_SZ 8

`define DDRMC5__PHY_RDEN4    32'h00000109
`define DDRMC5__PHY_RDEN4_SZ 8

`define DDRMC5__PHY_RDEN5    32'h0000010a
`define DDRMC5__PHY_RDEN5_SZ 8

`define DDRMC5__PHY_RDEN6    32'h0000010b
`define DDRMC5__PHY_RDEN6_SZ 8

`define DDRMC5__PHY_RDEN7    32'h0000010c
`define DDRMC5__PHY_RDEN7_SZ 8

`define DDRMC5__PHY_RDEN8    32'h0000010d
`define DDRMC5__PHY_RDEN8_SZ 8

`define DDRMC5__PHY_RDEN9    32'h0000010e
`define DDRMC5__PHY_RDEN9_SZ 8

`define DDRMC5__POWER_MANAGEMENT    32'h0000010f
`define DDRMC5__POWER_MANAGEMENT_SZ 28

`define DDRMC5__PRBS_MAX_LOOPS    32'h00000110
`define DDRMC5__PRBS_MAX_LOOPS_SZ 12

`define DDRMC5__PRBS_MAX_ROW_COL    32'h00000111
`define DDRMC5__PRBS_MAX_ROW_COL_SZ 25

`define DDRMC5__PRBS_SEED0    32'h00000112
`define DDRMC5__PRBS_SEED0_SZ 23

`define DDRMC5__PRBS_SEED1    32'h00000113
`define DDRMC5__PRBS_SEED1_SZ 23

`define DDRMC5__PRBS_SEED2    32'h00000114
`define DDRMC5__PRBS_SEED2_SZ 23

`define DDRMC5__PRBS_SEED3    32'h00000115
`define DDRMC5__PRBS_SEED3_SZ 23

`define DDRMC5__PRBS_SEED4    32'h00000116
`define DDRMC5__PRBS_SEED4_SZ 23

`define DDRMC5__PRBS_SEED5    32'h00000117
`define DDRMC5__PRBS_SEED5_SZ 23

`define DDRMC5__PRBS_SEED6    32'h00000118
`define DDRMC5__PRBS_SEED6_SZ 23

`define DDRMC5__PRBS_SEED7    32'h00000119
`define DDRMC5__PRBS_SEED7_SZ 23

`define DDRMC5__PRBS_SEED8    32'h0000011a
`define DDRMC5__PRBS_SEED8_SZ 23

`define DDRMC5__PRBS_TREF    32'h0000011b
`define DDRMC5__PRBS_TREF_SZ 24

`define DDRMC5__RAM_ERR_EN    32'h0000011c
`define DDRMC5__RAM_ERR_EN_SZ 7

`define DDRMC5__RAM_SETTING_RF2PHS    32'h0000011d
`define DDRMC5__RAM_SETTING_RF2PHS_SZ 8

`define DDRMC5__RAM_SETTING_RFSPHD    32'h0000011e
`define DDRMC5__RAM_SETTING_RFSPHD_SZ 7

`define DDRMC5__RAM_SETTING_SRSPHD    32'h0000011f
`define DDRMC5__RAM_SETTING_SRSPHD_SZ 7

`define DDRMC5__READ_DATA_EARLY_ID    32'h00000120
`define DDRMC5__READ_DATA_EARLY_ID_SZ 3

`define DDRMC5__REG_ADEC0    32'h00000121
`define DDRMC5__REG_ADEC0_SZ 20

`define DDRMC5__REG_ADEC1    32'h00000122
`define DDRMC5__REG_ADEC1_SZ 20

`define DDRMC5__REG_ADEC10    32'h00000123
`define DDRMC5__REG_ADEC10_SZ 30

`define DDRMC5__REG_ADEC11    32'h00000124
`define DDRMC5__REG_ADEC11_SZ 30

`define DDRMC5__REG_ADEC12    32'h00000125
`define DDRMC5__REG_ADEC12_SZ 30

`define DDRMC5__REG_ADEC13    32'h00000126
`define DDRMC5__REG_ADEC13_SZ 7

`define DDRMC5__REG_ADEC14    32'h00000127
`define DDRMC5__REG_ADEC14_SZ 29

`define DDRMC5__REG_ADEC15    32'h00000128
`define DDRMC5__REG_ADEC15_SZ 28

`define DDRMC5__REG_ADEC16    32'h00000129
`define DDRMC5__REG_ADEC16_SZ 32

`define DDRMC5__REG_ADEC2    32'h0000012a
`define DDRMC5__REG_ADEC2_SZ 21

`define DDRMC5__REG_ADEC3    32'h0000012b
`define DDRMC5__REG_ADEC3_SZ 20

`define DDRMC5__REG_ADEC4    32'h0000012c
`define DDRMC5__REG_ADEC4_SZ 12

`define DDRMC5__REG_ADEC5    32'h0000012d
`define DDRMC5__REG_ADEC5_SZ 24

`define DDRMC5__REG_ADEC6    32'h0000012e
`define DDRMC5__REG_ADEC6_SZ 30

`define DDRMC5__REG_ADEC7    32'h0000012f
`define DDRMC5__REG_ADEC7_SZ 30

`define DDRMC5__REG_ADEC8    32'h00000130
`define DDRMC5__REG_ADEC8_SZ 30

`define DDRMC5__REG_ADEC9    32'h00000131
`define DDRMC5__REG_ADEC9_SZ 30

`define DDRMC5__REG_ADEC_CHK0    32'h00000132
`define DDRMC5__REG_ADEC_CHK0_SZ 16

`define DDRMC5__REG_ADEC_CHK1    32'h00000133
`define DDRMC5__REG_ADEC_CHK1_SZ 32

`define DDRMC5__REG_ADEC_CHK2    32'h00000134
`define DDRMC5__REG_ADEC_CHK2_SZ 16

`define DDRMC5__REG_ADEC_CHK3    32'h00000135
`define DDRMC5__REG_ADEC_CHK3_SZ 32

`define DDRMC5__REG_ADEC_ILC    32'h00000136
`define DDRMC5__REG_ADEC_ILC_SZ 18

`define DDRMC5__REG_ADEC_MEMFILL0_HIGH    32'h00000137
`define DDRMC5__REG_ADEC_MEMFILL0_HIGH_SZ 32

`define DDRMC5__REG_ADEC_MEMFILL0_LOW    32'h00000138
`define DDRMC5__REG_ADEC_MEMFILL0_LOW_SZ 32

`define DDRMC5__REG_ADEC_MEMFILL1_HIGH    32'h00000139
`define DDRMC5__REG_ADEC_MEMFILL1_HIGH_SZ 32

`define DDRMC5__REG_ADEC_MEMFILL1_LOW    32'h0000013a
`define DDRMC5__REG_ADEC_MEMFILL1_LOW_SZ 32

`define DDRMC5__REG_AUTH_FAILURE    32'h0000013b
`define DDRMC5__REG_AUTH_FAILURE_SZ 16

`define DDRMC5__REG_CLKMON    32'h0000013c
`define DDRMC5__REG_CLKMON_SZ 6

`define DDRMC5__REG_CMDQ_BER_RATE_CTRL    32'h0000013d
`define DDRMC5__REG_CMDQ_BER_RATE_CTRL_SZ 22

`define DDRMC5__REG_CMDQ_BEW_RATE_CTRL    32'h0000013e
`define DDRMC5__REG_CMDQ_BEW_RATE_CTRL_SZ 22

`define DDRMC5__REG_CMDQ_ISR_RATE_CTRL    32'h0000013f
`define DDRMC5__REG_CMDQ_ISR_RATE_CTRL_SZ 22

`define DDRMC5__REG_CMDQ_ISW_RATE_CTRL    32'h00000140
`define DDRMC5__REG_CMDQ_ISW_RATE_CTRL_SZ 22

`define DDRMC5__REG_CMDQ_LLR_RATE_CTRL    32'h00000141
`define DDRMC5__REG_CMDQ_LLR_RATE_CTRL_SZ 22

`define DDRMC5__REG_COM_1    32'h00000142
`define DDRMC5__REG_COM_1_SZ 27

`define DDRMC5__REG_COM_2    32'h00000143
`define DDRMC5__REG_COM_2_SZ 27

`define DDRMC5__REG_COM_3    32'h00000144
`define DDRMC5__REG_COM_3_SZ 32

`define DDRMC5__REG_COM_6    32'h00000145
`define DDRMC5__REG_COM_6_SZ 14

`define DDRMC5__REG_CONFIG0    32'h00000146
`define DDRMC5__REG_CONFIG0_SZ 29

`define DDRMC5__REG_CONFIG1    32'h00000147
`define DDRMC5__REG_CONFIG1_SZ 3

`define DDRMC5__REG_CONFIG2    32'h00000148
`define DDRMC5__REG_CONFIG2_SZ 31

`define DDRMC5__REG_CONFIG3    32'h00000149
`define DDRMC5__REG_CONFIG3_SZ 32

`define DDRMC5__REG_CONFIG4    32'h0000014a
`define DDRMC5__REG_CONFIG4_SZ 24

`define DDRMC5__REG_CRP_ARB    32'h0000014b
`define DDRMC5__REG_CRP_ARB_SZ 16

`define DDRMC5__REG_CRYPTO_CTRL    32'h0000014c
`define DDRMC5__REG_CRYPTO_CTRL_SZ 32

`define DDRMC5__REG_CRYPTO_GCM_BM    32'h0000014d
`define DDRMC5__REG_CRYPTO_GCM_BM_SZ 8

`define DDRMC5__REG_CRYPTO_KEY_GEN    32'h0000014e
`define DDRMC5__REG_CRYPTO_KEY_GEN_SZ 24

`define DDRMC5__REG_CRYPTO_QOS    32'h0000014f
`define DDRMC5__REG_CRYPTO_QOS_SZ 32

`define DDRMC5__REG_CRYPTO_REKEY    32'h00000150
`define DDRMC5__REG_CRYPTO_REKEY_SZ 8

`define DDRMC5__REG_CRYPTO_XTS_BM    32'h00000151
`define DDRMC5__REG_CRYPTO_XTS_BM_SZ 8

`define DDRMC5__REG_DRAM_ARB    32'h00000152
`define DDRMC5__REG_DRAM_ARB_SZ 13

`define DDRMC5__REG_ERR_FATAL_EN    32'h00000153
`define DDRMC5__REG_ERR_FATAL_EN_SZ 26

`define DDRMC5__REG_ERR_NON_FATAL_EN    32'h00000154
`define DDRMC5__REG_ERR_NON_FATAL_EN_SZ 11

`define DDRMC5__REG_GCM0    32'h00000155
`define DDRMC5__REG_GCM0_SZ 32

`define DDRMC5__REG_GCM1    32'h00000156
`define DDRMC5__REG_GCM1_SZ 32

`define DDRMC5__REG_GCM10    32'h00000157
`define DDRMC5__REG_GCM10_SZ 32

`define DDRMC5__REG_GCM11    32'h00000158
`define DDRMC5__REG_GCM11_SZ 32

`define DDRMC5__REG_GCM12    32'h00000159
`define DDRMC5__REG_GCM12_SZ 32

`define DDRMC5__REG_GCM13    32'h0000015a
`define DDRMC5__REG_GCM13_SZ 32

`define DDRMC5__REG_GCM14    32'h0000015b
`define DDRMC5__REG_GCM14_SZ 32

`define DDRMC5__REG_GCM15    32'h0000015c
`define DDRMC5__REG_GCM15_SZ 32

`define DDRMC5__REG_GCM2    32'h0000015d
`define DDRMC5__REG_GCM2_SZ 32

`define DDRMC5__REG_GCM3    32'h0000015e
`define DDRMC5__REG_GCM3_SZ 32

`define DDRMC5__REG_GCM4    32'h0000015f
`define DDRMC5__REG_GCM4_SZ 32

`define DDRMC5__REG_GCM5    32'h00000160
`define DDRMC5__REG_GCM5_SZ 32

`define DDRMC5__REG_GCM6    32'h00000161
`define DDRMC5__REG_GCM6_SZ 32

`define DDRMC5__REG_GCM7    32'h00000162
`define DDRMC5__REG_GCM7_SZ 32

`define DDRMC5__REG_GCM8    32'h00000163
`define DDRMC5__REG_GCM8_SZ 32

`define DDRMC5__REG_GCM9    32'h00000164
`define DDRMC5__REG_GCM9_SZ 32

`define DDRMC5__REG_GCM_ILC    32'h00000165
`define DDRMC5__REG_GCM_ILC_SZ 32

`define DDRMC5__REG_KAT_ZEROIZE    32'h00000166
`define DDRMC5__REG_KAT_ZEROIZE_SZ 6

`define DDRMC5__REG_KEY_SCRUB    32'h00000167
`define DDRMC5__REG_KEY_SCRUB_SZ 6

`define DDRMC5__REG_META_C_SCRUB    32'h00000168
`define DDRMC5__REG_META_C_SCRUB_SZ 6

`define DDRMC5__REG_MRS_0    32'h00000169
`define DDRMC5__REG_MRS_0_SZ 28

`define DDRMC5__REG_MRS_1    32'h0000016a
`define DDRMC5__REG_MRS_1_SZ 32

`define DDRMC5__REG_MRS_2    32'h0000016b
`define DDRMC5__REG_MRS_2_SZ 4

`define DDRMC5__REG_MRS_7    32'h0000016c
`define DDRMC5__REG_MRS_7_SZ 12

`define DDRMC5__REG_NSU0_PORT    32'h0000016d
`define DDRMC5__REG_NSU0_PORT_SZ 12

`define DDRMC5__REG_NSU1_PORT    32'h0000016e
`define DDRMC5__REG_NSU1_PORT_SZ 12

`define DDRMC5__REG_NSU_0_EGR    32'h0000016f
`define DDRMC5__REG_NSU_0_EGR_SZ 30

`define DDRMC5__REG_NSU_0_ING    32'h00000170
`define DDRMC5__REG_NSU_0_ING_SZ 23

`define DDRMC5__REG_NSU_0_R_EGR    32'h00000171
`define DDRMC5__REG_NSU_0_R_EGR_SZ 28

`define DDRMC5__REG_NSU_0_W_EGR    32'h00000172
`define DDRMC5__REG_NSU_0_W_EGR_SZ 20

`define DDRMC5__REG_NSU_1_EGR    32'h00000173
`define DDRMC5__REG_NSU_1_EGR_SZ 30

`define DDRMC5__REG_NSU_1_ING    32'h00000174
`define DDRMC5__REG_NSU_1_ING_SZ 23

`define DDRMC5__REG_NSU_1_R_EGR    32'h00000175
`define DDRMC5__REG_NSU_1_R_EGR_SZ 28

`define DDRMC5__REG_NSU_1_W_EGR    32'h00000176
`define DDRMC5__REG_NSU_1_W_EGR_SZ 20

`define DDRMC5__REG_P0_BER_RATE_CTRL    32'h00000177
`define DDRMC5__REG_P0_BER_RATE_CTRL_SZ 22

`define DDRMC5__REG_P0_BEW_RATE_CTRL    32'h00000178
`define DDRMC5__REG_P0_BEW_RATE_CTRL_SZ 22

`define DDRMC5__REG_P0_ISR_RATE_CTRL    32'h00000179
`define DDRMC5__REG_P0_ISR_RATE_CTRL_SZ 22

`define DDRMC5__REG_P0_ISW_RATE_CTRL    32'h0000017a
`define DDRMC5__REG_P0_ISW_RATE_CTRL_SZ 22

`define DDRMC5__REG_P0_LLR_RATE_CTRL    32'h0000017b
`define DDRMC5__REG_P0_LLR_RATE_CTRL_SZ 22

`define DDRMC5__REG_P1_BER_RATE_CTRL    32'h0000017c
`define DDRMC5__REG_P1_BER_RATE_CTRL_SZ 22

`define DDRMC5__REG_P1_BEW_RATE_CTRL    32'h0000017d
`define DDRMC5__REG_P1_BEW_RATE_CTRL_SZ 22

`define DDRMC5__REG_P1_ISR_RATE_CTRL    32'h0000017e
`define DDRMC5__REG_P1_ISR_RATE_CTRL_SZ 22

`define DDRMC5__REG_P1_ISW_RATE_CTRL    32'h0000017f
`define DDRMC5__REG_P1_ISW_RATE_CTRL_SZ 22

`define DDRMC5__REG_P1_LLR_RATE_CTRL    32'h00000180
`define DDRMC5__REG_P1_LLR_RATE_CTRL_SZ 22

`define DDRMC5__REG_PINOUT    32'h00000181
`define DDRMC5__REG_PINOUT_SZ 19

`define DDRMC5__REG_PINOUT_ADDR_MUX_0    32'h00000182
`define DDRMC5__REG_PINOUT_ADDR_MUX_0_SZ 30

`define DDRMC5__REG_PINOUT_ADDR_MUX_1    32'h00000183
`define DDRMC5__REG_PINOUT_ADDR_MUX_1_SZ 30

`define DDRMC5__REG_PINOUT_ADDR_MUX_2    32'h00000184
`define DDRMC5__REG_PINOUT_ADDR_MUX_2_SZ 30

`define DDRMC5__REG_PT_CONFIG    32'h00000185
`define DDRMC5__REG_PT_CONFIG_SZ 20

`define DDRMC5__REG_QOS0    32'h00000186
`define DDRMC5__REG_QOS0_SZ 28

`define DDRMC5__REG_QOS1    32'h00000187
`define DDRMC5__REG_QOS1_SZ 30

`define DDRMC5__REG_QOS2    32'h00000188
`define DDRMC5__REG_QOS2_SZ 20

`define DDRMC5__REG_QOS_RATE_CTRL_SCALE    32'h00000189
`define DDRMC5__REG_QOS_RATE_CTRL_SCALE_SZ 25

`define DDRMC5__REG_QOS_TIMEOUT0    32'h0000018a
`define DDRMC5__REG_QOS_TIMEOUT0_SZ 25

`define DDRMC5__REG_QOS_TIMEOUT1    32'h0000018b
`define DDRMC5__REG_QOS_TIMEOUT1_SZ 32

`define DDRMC5__REG_QOS_TIMEOUT2    32'h0000018c
`define DDRMC5__REG_QOS_TIMEOUT2_SZ 8

`define DDRMC5__REG_RATE_CTRL_SCALE    32'h0000018d
`define DDRMC5__REG_RATE_CTRL_SCALE_SZ 25

`define DDRMC5__REG_RD_CONFIG    32'h0000018e
`define DDRMC5__REG_RD_CONFIG_SZ 6

`define DDRMC5__REG_RD_DRR_TKN_P0    32'h0000018f
`define DDRMC5__REG_RD_DRR_TKN_P0_SZ 24

`define DDRMC5__REG_RD_DRR_TKN_P1    32'h00000190
`define DDRMC5__REG_RD_DRR_TKN_P1_SZ 24

`define DDRMC5__REG_REF_0    32'h00000191
`define DDRMC5__REG_REF_0_SZ 3

`define DDRMC5__REG_REF_1    32'h00000192
`define DDRMC5__REG_REF_1_SZ 21

`define DDRMC5__REG_REF_2    32'h00000193
`define DDRMC5__REG_REF_2_SZ 3

`define DDRMC5__REG_REF_3    32'h00000194
`define DDRMC5__REG_REF_3_SZ 20

`define DDRMC5__REG_REF_4    32'h00000195
`define DDRMC5__REG_REF_4_SZ 2

`define DDRMC5__REG_REF_5    32'h00000196
`define DDRMC5__REG_REF_5_SZ 21

`define DDRMC5__REG_REF_6    32'h00000197
`define DDRMC5__REG_REF_6_SZ 1

`define DDRMC5__REG_REKEY_CTRL    32'h00000198
`define DDRMC5__REG_REKEY_CTRL_SZ 27

`define DDRMC5__REG_RETRY_0    32'h00000199
`define DDRMC5__REG_RETRY_0_SZ 29

`define DDRMC5__REG_RETRY_1    32'h0000019a
`define DDRMC5__REG_RETRY_1_SZ 30

`define DDRMC5__REG_RETRY_2    32'h0000019b
`define DDRMC5__REG_RETRY_2_SZ 29

`define DDRMC5__REG_RFM    32'h0000019c
`define DDRMC5__REG_RFM_SZ 29

`define DDRMC5__REG_RFM_1    32'h0000019d
`define DDRMC5__REG_RFM_1_SZ 11

`define DDRMC5__REG_SAFE_CONFIG0    32'h0000019e
`define DDRMC5__REG_SAFE_CONFIG0_SZ 26

`define DDRMC5__REG_SAFE_CONFIG1    32'h0000019f
`define DDRMC5__REG_SAFE_CONFIG1_SZ 32

`define DDRMC5__REG_SAFE_CONFIG10    32'h000001a0
`define DDRMC5__REG_SAFE_CONFIG10_SZ 32

`define DDRMC5__REG_SAFE_CONFIG11    32'h000001a1
`define DDRMC5__REG_SAFE_CONFIG11_SZ 28

`define DDRMC5__REG_SAFE_CONFIG12    32'h000001a2
`define DDRMC5__REG_SAFE_CONFIG12_SZ 24

`define DDRMC5__REG_SAFE_CONFIG13    32'h000001a3
`define DDRMC5__REG_SAFE_CONFIG13_SZ 24

`define DDRMC5__REG_SAFE_CONFIG14    32'h000001a4
`define DDRMC5__REG_SAFE_CONFIG14_SZ 32

`define DDRMC5__REG_SAFE_CONFIG15    32'h000001a5
`define DDRMC5__REG_SAFE_CONFIG15_SZ 32

`define DDRMC5__REG_SAFE_CONFIG2    32'h000001a6
`define DDRMC5__REG_SAFE_CONFIG2_SZ 30

`define DDRMC5__REG_SAFE_CONFIG3    32'h000001a7
`define DDRMC5__REG_SAFE_CONFIG3_SZ 32

`define DDRMC5__REG_SAFE_CONFIG4    32'h000001a8
`define DDRMC5__REG_SAFE_CONFIG4_SZ 29

`define DDRMC5__REG_SAFE_CONFIG5    32'h000001a9
`define DDRMC5__REG_SAFE_CONFIG5_SZ 32

`define DDRMC5__REG_SAFE_CONFIG6    32'h000001aa
`define DDRMC5__REG_SAFE_CONFIG6_SZ 31

`define DDRMC5__REG_SAFE_CONFIG7    32'h000001ab
`define DDRMC5__REG_SAFE_CONFIG7_SZ 32

`define DDRMC5__REG_SAFE_CONFIG8    32'h000001ac
`define DDRMC5__REG_SAFE_CONFIG8_SZ 32

`define DDRMC5__REG_SAFE_CONFIG9    32'h000001ad
`define DDRMC5__REG_SAFE_CONFIG9_SZ 32

`define DDRMC5__REG_SAFE_MUX    32'h000001ae
`define DDRMC5__REG_SAFE_MUX_SZ 2

`define DDRMC5__REG_SCRUB_ADDR_RANGE_HI    32'h000001af
`define DDRMC5__REG_SCRUB_ADDR_RANGE_HI_SZ 4

`define DDRMC5__REG_SCRUB_ADDR_RANGE_LO    32'h000001b0
`define DDRMC5__REG_SCRUB_ADDR_RANGE_LO_SZ 32

`define DDRMC5__REG_SCRUB_BASE_ADDR_HI    32'h000001b1
`define DDRMC5__REG_SCRUB_BASE_ADDR_HI_SZ 16

`define DDRMC5__REG_SCRUB_BASE_ADDR_LO    32'h000001b2
`define DDRMC5__REG_SCRUB_BASE_ADDR_LO_SZ 32

`define DDRMC5__REG_SCRUB_CONFIG    32'h000001b3
`define DDRMC5__REG_SCRUB_CONFIG_SZ 5

`define DDRMC5__REG_SCRUB_DEBUG_MODE    32'h000001b4
`define DDRMC5__REG_SCRUB_DEBUG_MODE_SZ 2

`define DDRMC5__REG_SCRUB_INTVL    32'h000001b5
`define DDRMC5__REG_SCRUB_INTVL_SZ 24

`define DDRMC5__REG_SCRUB_OTF    32'h000001b6
`define DDRMC5__REG_SCRUB_OTF_SZ 2

`define DDRMC5__REG_SCRUB_PER_RD    32'h000001b7
`define DDRMC5__REG_SCRUB_PER_RD_SZ 32

`define DDRMC5__REG_SCRUB_TAP    32'h000001b8
`define DDRMC5__REG_SCRUB_TAP_SZ 24

`define DDRMC5__REG_SCRUB_TO    32'h000001b9
`define DDRMC5__REG_SCRUB_TO_SZ 32

`define DDRMC5__REG_SCRUB_WAIT    32'h000001ba
`define DDRMC5__REG_SCRUB_WAIT_SZ 8

`define DDRMC5__REG_SND_AUTH_SCRUB    32'h000001bb
`define DDRMC5__REG_SND_AUTH_SCRUB_SZ 6

`define DDRMC5__REG_TIMER_FIFO    32'h000001bc
`define DDRMC5__REG_TIMER_FIFO_SZ 6

`define DDRMC5__REG_TXN_CONFIG    32'h000001bd
`define DDRMC5__REG_TXN_CONFIG_SZ 28

`define DDRMC5__REG_TXN_CONFIG_1    32'h000001be
`define DDRMC5__REG_TXN_CONFIG_1_SZ 32

`define DDRMC5__REG_TXN_CONFIG_2    32'h000001bf
`define DDRMC5__REG_TXN_CONFIG_2_SZ 7

`define DDRMC5__REG_TXN_CONFIG_3    32'h000001c0
`define DDRMC5__REG_TXN_CONFIG_3_SZ 16

`define DDRMC5__REG_WR_CONFIG    32'h000001c1
`define DDRMC5__REG_WR_CONFIG_SZ 32

`define DDRMC5__REG_WR_DRR_TKN_P0    32'h000001c2
`define DDRMC5__REG_WR_DRR_TKN_P0_SZ 16

`define DDRMC5__REG_WR_DRR_TKN_P1    32'h000001c3
`define DDRMC5__REG_WR_DRR_TKN_P1_SZ 16

`define DDRMC5__TRSS_TIMEOUT    32'h000001c4
`define DDRMC5__TRSS_TIMEOUT_SZ 6

`define DDRMC5__TXNQ_ENTRY_COUNT_MODE    32'h000001c5
`define DDRMC5__TXNQ_ENTRY_COUNT_MODE_SZ 14

`define DDRMC5__TXNQ_RD_PRIORITY    32'h000001c6
`define DDRMC5__TXNQ_RD_PRIORITY_SZ 26

`define DDRMC5__TXNQ_WR_PRIORITY    32'h000001c7
`define DDRMC5__TXNQ_WR_PRIORITY_SZ 25

`define DDRMC5__UB_CLK_MUX    32'h000001c8
`define DDRMC5__UB_CLK_MUX_SZ 2

`define DDRMC5__X5PHYIO_STARTUP    32'h000001c9
`define DDRMC5__X5PHYIO_STARTUP_SZ 8

`define DDRMC5__XMPU_CONFIG0    32'h000001ca
`define DDRMC5__XMPU_CONFIG0_SZ 5

`define DDRMC5__XMPU_CONFIG1    32'h000001cb
`define DDRMC5__XMPU_CONFIG1_SZ 5

`define DDRMC5__XMPU_CONFIG10    32'h000001cc
`define DDRMC5__XMPU_CONFIG10_SZ 5

`define DDRMC5__XMPU_CONFIG11    32'h000001cd
`define DDRMC5__XMPU_CONFIG11_SZ 5

`define DDRMC5__XMPU_CONFIG12    32'h000001ce
`define DDRMC5__XMPU_CONFIG12_SZ 5

`define DDRMC5__XMPU_CONFIG13    32'h000001cf
`define DDRMC5__XMPU_CONFIG13_SZ 5

`define DDRMC5__XMPU_CONFIG14    32'h000001d0
`define DDRMC5__XMPU_CONFIG14_SZ 5

`define DDRMC5__XMPU_CONFIG15    32'h000001d1
`define DDRMC5__XMPU_CONFIG15_SZ 5

`define DDRMC5__XMPU_CONFIG2    32'h000001d2
`define DDRMC5__XMPU_CONFIG2_SZ 5

`define DDRMC5__XMPU_CONFIG3    32'h000001d3
`define DDRMC5__XMPU_CONFIG3_SZ 5

`define DDRMC5__XMPU_CONFIG4    32'h000001d4
`define DDRMC5__XMPU_CONFIG4_SZ 5

`define DDRMC5__XMPU_CONFIG5    32'h000001d5
`define DDRMC5__XMPU_CONFIG5_SZ 5

`define DDRMC5__XMPU_CONFIG6    32'h000001d6
`define DDRMC5__XMPU_CONFIG6_SZ 5

`define DDRMC5__XMPU_CONFIG7    32'h000001d7
`define DDRMC5__XMPU_CONFIG7_SZ 5

`define DDRMC5__XMPU_CONFIG8    32'h000001d8
`define DDRMC5__XMPU_CONFIG8_SZ 5

`define DDRMC5__XMPU_CONFIG9    32'h000001d9
`define DDRMC5__XMPU_CONFIG9_SZ 5

`define DDRMC5__XMPU_CRPTO_CFG0_0    32'h000001da
`define DDRMC5__XMPU_CRPTO_CFG0_0_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_1    32'h000001db
`define DDRMC5__XMPU_CRPTO_CFG0_1_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_10    32'h000001dc
`define DDRMC5__XMPU_CRPTO_CFG0_10_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_11    32'h000001dd
`define DDRMC5__XMPU_CRPTO_CFG0_11_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_12    32'h000001de
`define DDRMC5__XMPU_CRPTO_CFG0_12_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_13    32'h000001df
`define DDRMC5__XMPU_CRPTO_CFG0_13_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_14    32'h000001e0
`define DDRMC5__XMPU_CRPTO_CFG0_14_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_15    32'h000001e1
`define DDRMC5__XMPU_CRPTO_CFG0_15_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_2    32'h000001e2
`define DDRMC5__XMPU_CRPTO_CFG0_2_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_3    32'h000001e3
`define DDRMC5__XMPU_CRPTO_CFG0_3_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_4    32'h000001e4
`define DDRMC5__XMPU_CRPTO_CFG0_4_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_5    32'h000001e5
`define DDRMC5__XMPU_CRPTO_CFG0_5_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_6    32'h000001e6
`define DDRMC5__XMPU_CRPTO_CFG0_6_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_7    32'h000001e7
`define DDRMC5__XMPU_CRPTO_CFG0_7_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_8    32'h000001e8
`define DDRMC5__XMPU_CRPTO_CFG0_8_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG0_9    32'h000001e9
`define DDRMC5__XMPU_CRPTO_CFG0_9_SZ 8

`define DDRMC5__XMPU_CRPTO_CFG1_0    32'h000001ea
`define DDRMC5__XMPU_CRPTO_CFG1_0_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_1    32'h000001eb
`define DDRMC5__XMPU_CRPTO_CFG1_1_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_10    32'h000001ec
`define DDRMC5__XMPU_CRPTO_CFG1_10_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_11    32'h000001ed
`define DDRMC5__XMPU_CRPTO_CFG1_11_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_12    32'h000001ee
`define DDRMC5__XMPU_CRPTO_CFG1_12_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_13    32'h000001ef
`define DDRMC5__XMPU_CRPTO_CFG1_13_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_14    32'h000001f0
`define DDRMC5__XMPU_CRPTO_CFG1_14_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_15    32'h000001f1
`define DDRMC5__XMPU_CRPTO_CFG1_15_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_2    32'h000001f2
`define DDRMC5__XMPU_CRPTO_CFG1_2_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_3    32'h000001f3
`define DDRMC5__XMPU_CRPTO_CFG1_3_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_4    32'h000001f4
`define DDRMC5__XMPU_CRPTO_CFG1_4_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_5    32'h000001f5
`define DDRMC5__XMPU_CRPTO_CFG1_5_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_6    32'h000001f6
`define DDRMC5__XMPU_CRPTO_CFG1_6_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_7    32'h000001f7
`define DDRMC5__XMPU_CRPTO_CFG1_7_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_8    32'h000001f8
`define DDRMC5__XMPU_CRPTO_CFG1_8_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG1_9    32'h000001f9
`define DDRMC5__XMPU_CRPTO_CFG1_9_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_0    32'h000001fa
`define DDRMC5__XMPU_CRPTO_CFG2_0_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_1    32'h000001fb
`define DDRMC5__XMPU_CRPTO_CFG2_1_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_10    32'h000001fc
`define DDRMC5__XMPU_CRPTO_CFG2_10_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_11    32'h000001fd
`define DDRMC5__XMPU_CRPTO_CFG2_11_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_12    32'h000001fe
`define DDRMC5__XMPU_CRPTO_CFG2_12_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_13    32'h000001ff
`define DDRMC5__XMPU_CRPTO_CFG2_13_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_14    32'h00000200
`define DDRMC5__XMPU_CRPTO_CFG2_14_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_15    32'h00000201
`define DDRMC5__XMPU_CRPTO_CFG2_15_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_2    32'h00000202
`define DDRMC5__XMPU_CRPTO_CFG2_2_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_3    32'h00000203
`define DDRMC5__XMPU_CRPTO_CFG2_3_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_4    32'h00000204
`define DDRMC5__XMPU_CRPTO_CFG2_4_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_5    32'h00000205
`define DDRMC5__XMPU_CRPTO_CFG2_5_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_6    32'h00000206
`define DDRMC5__XMPU_CRPTO_CFG2_6_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_7    32'h00000207
`define DDRMC5__XMPU_CRPTO_CFG2_7_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_8    32'h00000208
`define DDRMC5__XMPU_CRPTO_CFG2_8_SZ 28

`define DDRMC5__XMPU_CRPTO_CFG2_9    32'h00000209
`define DDRMC5__XMPU_CRPTO_CFG2_9_SZ 28

`define DDRMC5__XMPU_CTRL    32'h0000020a
`define DDRMC5__XMPU_CTRL_SZ 7

`define DDRMC5__XMPU_END_HI0    32'h0000020b
`define DDRMC5__XMPU_END_HI0_SZ 16

`define DDRMC5__XMPU_END_HI1    32'h0000020c
`define DDRMC5__XMPU_END_HI1_SZ 16

`define DDRMC5__XMPU_END_HI10    32'h0000020d
`define DDRMC5__XMPU_END_HI10_SZ 16

`define DDRMC5__XMPU_END_HI11    32'h0000020e
`define DDRMC5__XMPU_END_HI11_SZ 16

`define DDRMC5__XMPU_END_HI12    32'h0000020f
`define DDRMC5__XMPU_END_HI12_SZ 16

`define DDRMC5__XMPU_END_HI13    32'h00000210
`define DDRMC5__XMPU_END_HI13_SZ 16

`define DDRMC5__XMPU_END_HI14    32'h00000211
`define DDRMC5__XMPU_END_HI14_SZ 16

`define DDRMC5__XMPU_END_HI15    32'h00000212
`define DDRMC5__XMPU_END_HI15_SZ 16

`define DDRMC5__XMPU_END_HI2    32'h00000213
`define DDRMC5__XMPU_END_HI2_SZ 16

`define DDRMC5__XMPU_END_HI3    32'h00000214
`define DDRMC5__XMPU_END_HI3_SZ 16

`define DDRMC5__XMPU_END_HI4    32'h00000215
`define DDRMC5__XMPU_END_HI4_SZ 16

`define DDRMC5__XMPU_END_HI5    32'h00000216
`define DDRMC5__XMPU_END_HI5_SZ 16

`define DDRMC5__XMPU_END_HI6    32'h00000217
`define DDRMC5__XMPU_END_HI6_SZ 16

`define DDRMC5__XMPU_END_HI7    32'h00000218
`define DDRMC5__XMPU_END_HI7_SZ 16

`define DDRMC5__XMPU_END_HI8    32'h00000219
`define DDRMC5__XMPU_END_HI8_SZ 16

`define DDRMC5__XMPU_END_HI9    32'h0000021a
`define DDRMC5__XMPU_END_HI9_SZ 16

`define DDRMC5__XMPU_END_LO0    32'h0000021b
`define DDRMC5__XMPU_END_LO0_SZ 32

`define DDRMC5__XMPU_END_LO1    32'h0000021c
`define DDRMC5__XMPU_END_LO1_SZ 32

`define DDRMC5__XMPU_END_LO10    32'h0000021d
`define DDRMC5__XMPU_END_LO10_SZ 32

`define DDRMC5__XMPU_END_LO11    32'h0000021e
`define DDRMC5__XMPU_END_LO11_SZ 32

`define DDRMC5__XMPU_END_LO12    32'h0000021f
`define DDRMC5__XMPU_END_LO12_SZ 32

`define DDRMC5__XMPU_END_LO13    32'h00000220
`define DDRMC5__XMPU_END_LO13_SZ 32

`define DDRMC5__XMPU_END_LO14    32'h00000221
`define DDRMC5__XMPU_END_LO14_SZ 32

`define DDRMC5__XMPU_END_LO15    32'h00000222
`define DDRMC5__XMPU_END_LO15_SZ 32

`define DDRMC5__XMPU_END_LO2    32'h00000223
`define DDRMC5__XMPU_END_LO2_SZ 32

`define DDRMC5__XMPU_END_LO3    32'h00000224
`define DDRMC5__XMPU_END_LO3_SZ 32

`define DDRMC5__XMPU_END_LO4    32'h00000225
`define DDRMC5__XMPU_END_LO4_SZ 32

`define DDRMC5__XMPU_END_LO5    32'h00000226
`define DDRMC5__XMPU_END_LO5_SZ 32

`define DDRMC5__XMPU_END_LO6    32'h00000227
`define DDRMC5__XMPU_END_LO6_SZ 32

`define DDRMC5__XMPU_END_LO7    32'h00000228
`define DDRMC5__XMPU_END_LO7_SZ 32

`define DDRMC5__XMPU_END_LO8    32'h00000229
`define DDRMC5__XMPU_END_LO8_SZ 32

`define DDRMC5__XMPU_END_LO9    32'h0000022a
`define DDRMC5__XMPU_END_LO9_SZ 32

`define DDRMC5__XMPU_MASTER0    32'h0000022b
`define DDRMC5__XMPU_MASTER0_SZ 26

`define DDRMC5__XMPU_MASTER1    32'h0000022c
`define DDRMC5__XMPU_MASTER1_SZ 26

`define DDRMC5__XMPU_MASTER10    32'h0000022d
`define DDRMC5__XMPU_MASTER10_SZ 26

`define DDRMC5__XMPU_MASTER11    32'h0000022e
`define DDRMC5__XMPU_MASTER11_SZ 26

`define DDRMC5__XMPU_MASTER12    32'h0000022f
`define DDRMC5__XMPU_MASTER12_SZ 26

`define DDRMC5__XMPU_MASTER13    32'h00000230
`define DDRMC5__XMPU_MASTER13_SZ 26

`define DDRMC5__XMPU_MASTER14    32'h00000231
`define DDRMC5__XMPU_MASTER14_SZ 26

`define DDRMC5__XMPU_MASTER15    32'h00000232
`define DDRMC5__XMPU_MASTER15_SZ 26

`define DDRMC5__XMPU_MASTER2    32'h00000233
`define DDRMC5__XMPU_MASTER2_SZ 26

`define DDRMC5__XMPU_MASTER3    32'h00000234
`define DDRMC5__XMPU_MASTER3_SZ 26

`define DDRMC5__XMPU_MASTER4    32'h00000235
`define DDRMC5__XMPU_MASTER4_SZ 26

`define DDRMC5__XMPU_MASTER5    32'h00000236
`define DDRMC5__XMPU_MASTER5_SZ 26

`define DDRMC5__XMPU_MASTER6    32'h00000237
`define DDRMC5__XMPU_MASTER6_SZ 26

`define DDRMC5__XMPU_MASTER7    32'h00000238
`define DDRMC5__XMPU_MASTER7_SZ 26

`define DDRMC5__XMPU_MASTER8    32'h00000239
`define DDRMC5__XMPU_MASTER8_SZ 26

`define DDRMC5__XMPU_MASTER9    32'h0000023a
`define DDRMC5__XMPU_MASTER9_SZ 26

`define DDRMC5__XMPU_START_HI0    32'h0000023b
`define DDRMC5__XMPU_START_HI0_SZ 16

`define DDRMC5__XMPU_START_HI1    32'h0000023c
`define DDRMC5__XMPU_START_HI1_SZ 16

`define DDRMC5__XMPU_START_HI10    32'h0000023d
`define DDRMC5__XMPU_START_HI10_SZ 16

`define DDRMC5__XMPU_START_HI11    32'h0000023e
`define DDRMC5__XMPU_START_HI11_SZ 16

`define DDRMC5__XMPU_START_HI12    32'h0000023f
`define DDRMC5__XMPU_START_HI12_SZ 16

`define DDRMC5__XMPU_START_HI13    32'h00000240
`define DDRMC5__XMPU_START_HI13_SZ 16

`define DDRMC5__XMPU_START_HI14    32'h00000241
`define DDRMC5__XMPU_START_HI14_SZ 16

`define DDRMC5__XMPU_START_HI15    32'h00000242
`define DDRMC5__XMPU_START_HI15_SZ 16

`define DDRMC5__XMPU_START_HI2    32'h00000243
`define DDRMC5__XMPU_START_HI2_SZ 16

`define DDRMC5__XMPU_START_HI3    32'h00000244
`define DDRMC5__XMPU_START_HI3_SZ 16

`define DDRMC5__XMPU_START_HI4    32'h00000245
`define DDRMC5__XMPU_START_HI4_SZ 16

`define DDRMC5__XMPU_START_HI5    32'h00000246
`define DDRMC5__XMPU_START_HI5_SZ 16

`define DDRMC5__XMPU_START_HI6    32'h00000247
`define DDRMC5__XMPU_START_HI6_SZ 16

`define DDRMC5__XMPU_START_HI7    32'h00000248
`define DDRMC5__XMPU_START_HI7_SZ 16

`define DDRMC5__XMPU_START_HI8    32'h00000249
`define DDRMC5__XMPU_START_HI8_SZ 16

`define DDRMC5__XMPU_START_HI9    32'h0000024a
`define DDRMC5__XMPU_START_HI9_SZ 16

`define DDRMC5__XMPU_START_LO0    32'h0000024b
`define DDRMC5__XMPU_START_LO0_SZ 32

`define DDRMC5__XMPU_START_LO1    32'h0000024c
`define DDRMC5__XMPU_START_LO1_SZ 32

`define DDRMC5__XMPU_START_LO10    32'h0000024d
`define DDRMC5__XMPU_START_LO10_SZ 32

`define DDRMC5__XMPU_START_LO11    32'h0000024e
`define DDRMC5__XMPU_START_LO11_SZ 32

`define DDRMC5__XMPU_START_LO12    32'h0000024f
`define DDRMC5__XMPU_START_LO12_SZ 32

`define DDRMC5__XMPU_START_LO13    32'h00000250
`define DDRMC5__XMPU_START_LO13_SZ 32

`define DDRMC5__XMPU_START_LO14    32'h00000251
`define DDRMC5__XMPU_START_LO14_SZ 32

`define DDRMC5__XMPU_START_LO15    32'h00000252
`define DDRMC5__XMPU_START_LO15_SZ 32

`define DDRMC5__XMPU_START_LO2    32'h00000253
`define DDRMC5__XMPU_START_LO2_SZ 32

`define DDRMC5__XMPU_START_LO3    32'h00000254
`define DDRMC5__XMPU_START_LO3_SZ 32

`define DDRMC5__XMPU_START_LO4    32'h00000255
`define DDRMC5__XMPU_START_LO4_SZ 32

`define DDRMC5__XMPU_START_LO5    32'h00000256
`define DDRMC5__XMPU_START_LO5_SZ 32

`define DDRMC5__XMPU_START_LO6    32'h00000257
`define DDRMC5__XMPU_START_LO6_SZ 32

`define DDRMC5__XMPU_START_LO7    32'h00000258
`define DDRMC5__XMPU_START_LO7_SZ 32

`define DDRMC5__XMPU_START_LO8    32'h00000259
`define DDRMC5__XMPU_START_LO8_SZ 32

`define DDRMC5__XMPU_START_LO9    32'h0000025a
`define DDRMC5__XMPU_START_LO9_SZ 32

`define DDRMC5__XPI_ADDR_CFG    32'h0000025b
`define DDRMC5__XPI_ADDR_CFG_SZ 5

`define DDRMC5__XPI_DQS_T_CNTRL    32'h0000025c
`define DDRMC5__XPI_DQS_T_CNTRL_SZ 24

`define DDRMC5__XPI_DQS_T_CNTRL_PREAMBLE0    32'h0000025d
`define DDRMC5__XPI_DQS_T_CNTRL_PREAMBLE0_SZ 32

`define DDRMC5__XPI_DQS_T_CNTRL_PREAMBLE1    32'h0000025e
`define DDRMC5__XPI_DQS_T_CNTRL_PREAMBLE1_SZ 32

`define DDRMC5__XPI_IBUF_DIS_OR_HS_RX_DIS    32'h0000025f
`define DDRMC5__XPI_IBUF_DIS_OR_HS_RX_DIS_SZ 7

`define DDRMC5__XPI_MAP_AC_TIE_OFF    32'h00000260
`define DDRMC5__XPI_MAP_AC_TIE_OFF_SZ 5

`define DDRMC5__XPI_MAP_CS_OVERRIDE_CFG    32'h00000261
`define DDRMC5__XPI_MAP_CS_OVERRIDE_CFG_SZ 2

`define DDRMC5__XPI_MAP_PD_EN    32'h00000262
`define DDRMC5__XPI_MAP_PD_EN_SZ 12

`define DDRMC5__XPI_MRS_CONFIG    32'h00000263
`define DDRMC5__XPI_MRS_CONFIG_SZ 16

`define DDRMC5__XPI_NON_TARGET_ODT    32'h00000264
`define DDRMC5__XPI_NON_TARGET_ODT_SZ 1

`define DDRMC5__XPI_NON_TARGET_ODT_CFG_READ    32'h00000265
`define DDRMC5__XPI_NON_TARGET_ODT_CFG_READ_SZ 16

`define DDRMC5__XPI_NON_TARGET_ODT_CFG_WRITE    32'h00000266
`define DDRMC5__XPI_NON_TARGET_ODT_CFG_WRITE_SZ 16

`define DDRMC5__XPI_OE_ALL_NIB    32'h00000267
`define DDRMC5__XPI_OE_ALL_NIB_SZ 11

`define DDRMC5__XPI_OE_CNTRL    32'h00000268
`define DDRMC5__XPI_OE_CNTRL_SZ 31

`define DDRMC5__XPI_OE_CNTRL2    32'h00000269
`define DDRMC5__XPI_OE_CNTRL2_SZ 4

`define DDRMC5__XPI_OE_CNTRL_PREAMBLE    32'h0000026a
`define DDRMC5__XPI_OE_CNTRL_PREAMBLE_SZ 32

`define DDRMC5__XPI_PMI_CONFIG    32'h0000026b
`define DDRMC5__XPI_PMI_CONFIG_SZ 2

`define DDRMC5__XPI_READ_DBI    32'h0000026c
`define DDRMC5__XPI_READ_DBI_SZ 1

`define DDRMC5__XPI_READ_NIB_ENABLE    32'h0000026d
`define DDRMC5__XPI_READ_NIB_ENABLE_SZ 10

`define DDRMC5__XPI_READ_OFFSET    32'h0000026e
`define DDRMC5__XPI_READ_OFFSET_SZ 15

`define DDRMC5__XPI_WRDATA_ALL_NIB    32'h0000026f
`define DDRMC5__XPI_WRDATA_ALL_NIB_SZ 15

`define DDRMC5__XPI_WRITE_DM_DBI    32'h00000270
`define DDRMC5__XPI_WRITE_DM_DBI_SZ 5

`define DDRMC5__XPI_WRITE_NIB_ENABLE    32'h00000271
`define DDRMC5__XPI_WRITE_NIB_ENABLE_SZ 10

`endif  // B_DDRMC5_DEFINES_VH