`include "B_IBUF_INTERMDISABLE_defines.vh"

reg [`IBUF_INTERMDISABLE_DATA_SZ-1:0] ATTR [0:`IBUF_INTERMDISABLE_ADDR_N-1];
reg [`IBUF_INTERMDISABLE__IBUF_LOW_PWR_SZ:1] IBUF_LOW_PWR_REG = IBUF_LOW_PWR;
reg [`IBUF_INTERMDISABLE__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IBUF_INTERMDISABLE__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`IBUF_INTERMDISABLE__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IBUF_INTERMDISABLE__IBUF_LOW_PWR] = IBUF_LOW_PWR;
  ATTR[`IBUF_INTERMDISABLE__IOSTANDARD] = IOSTANDARD;
  ATTR[`IBUF_INTERMDISABLE__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`IBUF_INTERMDISABLE__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  IBUF_LOW_PWR_REG = ATTR[`IBUF_INTERMDISABLE__IBUF_LOW_PWR];
  IOSTANDARD_REG = ATTR[`IBUF_INTERMDISABLE__IOSTANDARD];
  SIM_DEVICE_REG = ATTR[`IBUF_INTERMDISABLE__SIM_DEVICE];
  USE_IBUFDISABLE_REG = ATTR[`IBUF_INTERMDISABLE__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IBUF_INTERMDISABLE_ADDR_SZ-1:0] addr;
  input  [`IBUF_INTERMDISABLE_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IBUF_INTERMDISABLE_DATA_SZ-1:0] read_attr;
  input  [`IBUF_INTERMDISABLE_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
