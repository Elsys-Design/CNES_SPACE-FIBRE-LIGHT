-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 02/07/2025
--
-- Description : This module manages the reset of the Spacefibre hssl ip
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_init_hssl is
   port (
      RST_N                            : in  std_logic;    --! global reset
      CLK                              : in  std_logic;    --! Clock generated by HSSL IP
      -- PLSH interface
      PLL_PMA_PWR_UP_PLIH              : out std_logic;
      TX_DRIVER_PWRDWN_N_PLIH          : out std_logic;
      PLL_PMA_RST_N_PLIH               : out std_logic;
      PLL_PMA_LOCK_ANALOG_HSSL         : in  std_logic;
      TX_RST_N_PLIH                    : out std_logic;
      TX_BUSY_HSSL                     : in  std_logic;
      RX_PMA_PWR_UP_PLIH               : out std_logic;
      RX_PMA_RST_N_PLIH                : out std_logic;
      RX_PMA_LL_SLOW_LOCKED_HSSL       : in  std_logic;
      RX_RST_N_PLIH                    : out std_logic;
      RX_BUSY_HSSL                     : in  std_logic;
      -- Output
      HSSL_RESET_DONE_PLIH             : out std_logic
   );
end ppl_init_hssl;

architecture rtl of ppl_init_hssl is
---------------------------------------------------------
-----                   Type declaration            -----
---------------------------------------------------------
  type ppl_pma_pll_fsm is (
    PMA_PLL_POWER_UP_ST,
    TX_POWER_UP_ST,
    PMA_PLL_RST_PULSE_ST,
    PMA_PLL_LOCK_ST
  );

  type ppl_rx_pma_pll_fsm is (
    IDLE_ST,
    RX_PMA_POWER_UP_ST,
    RX_PMA_PLL_PULSE_ST,
    RX_PMA_LOCK_ST,
    RX_RST_PULSE_ST,
    RX_STARTED_ST
  );

  type ppl_tx_pcs_fsm is (
    IDLE_ST,
    TX_PULSE_ST,
    TX_STARTED_ST
  );
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
  signal current_state_pll_pma      : ppl_pma_pll_fsm;
  signal current_state_rx_pll_pma   : ppl_rx_pma_pll_fsm;
  signal current_state_tx_pcs       : ppl_tx_pcs_fsm;
  signal pma_pll_seq_end            : std_logic;
  signal rx_pll_pma_started         : std_logic;
  signal tx_pcs_started             : std_logic;

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_pma_pll
-- Description: Manages the PMA PLL reset of the SpaceFibre
--              HSSL IP
---------------------------------------------------------
p_pma_pll: process(CLK, RST_N)
begin
  if RST_N ='0' then
    current_state_pll_pma   <= PMA_PLL_POWER_UP_ST;
    PLL_PMA_PWR_UP_PLIH     <= '0';
    TX_DRIVER_PWRDWN_N_PLIH <= '0';
    PLL_PMA_RST_N_PLIH      <= '0';
    pma_pll_seq_end         <= '0';
  elsif rising_edge(CLK)  then
    case current_state_pll_pma is
      when PMA_PLL_POWER_UP_ST =>
                                    PLL_PMA_PWR_UP_PLIH   <= '1'; -- PMA PLL power up
                                    current_state_pll_pma <= TX_POWER_UP_ST;
      when TX_POWER_UP_ST =>
                                    TX_DRIVER_PWRDWN_N_PLIH <= '1'; -- TX driver power up
                                    current_state_pll_pma   <= PMA_PLL_RST_PULSE_ST;
      when PMA_PLL_RST_PULSE_ST =>
                                    PLL_PMA_RST_N_PLIH      <= '1'; -- PMA PLL rst pulse
                                    current_state_pll_pma <= PMA_PLL_LOCK_ST;
      when PMA_PLL_LOCK_ST =>
                                    if PLL_PMA_LOCK_ANALOG_HSSL ='1' then -- PMA PLL is locked
                                      pma_pll_seq_end <= '1';
                                    end if;
      when others =>
                                    current_state_pll_pma <= PMA_PLL_POWER_UP_ST;
    end case;
  end if;
end process p_pma_pll;

---------------------------------------------------------
-- Process: p_rx_pma_pll
-- Description: Manages the RX PMA PLL and RX PCS reset
--              of the SpaceFibre HSSL IP
---------------------------------------------------------
p_rx_pma_pll: process(CLK, RST_N)
begin
  if RST_N ='0' then
    current_state_rx_pll_pma <= IDLE_ST;
    RX_PMA_PWR_UP_PLIH       <= '0';
    RX_PMA_RST_N_PLIH        <= '0';
    RX_RST_N_PLIH            <= '0';
    rx_pll_pma_started       <= '0';
  elsif rising_edge(CLK)  then
    rx_pll_pma_started <= '0';
    case current_state_rx_pll_pma is
      when IDLE_ST =>
                                    if pma_pll_seq_end = '1' then -- PMA PLL is locked
                                      current_state_rx_pll_pma <= RX_PMA_POWER_UP_ST;
                                    end if;
      when RX_PMA_POWER_UP_ST =>
                                    RX_PMA_PWR_UP_PLIH         <= '1'; -- RX PMA power up
                                    current_state_rx_pll_pma   <= RX_PMA_PLL_PULSE_ST;
      when RX_PMA_PLL_PULSE_ST =>
                                    RX_PMA_RST_N_PLIH        <= '1';-- RX PMA PLL rst pulse
                                    current_state_rx_pll_pma <= RX_PMA_LOCK_ST;
      when RX_PMA_LOCK_ST =>
                                    if RX_PMA_LL_SLOW_LOCKED_HSSL ='1' then -- RX PMA PLL is locked
                                      current_state_rx_pll_pma <= RX_RST_PULSE_ST;
                                    end if;
      when RX_RST_PULSE_ST =>
                                    RX_RST_N_PLIH            <= '1'; -- RX PCS rst pulse
                                    current_state_rx_pll_pma <= RX_STARTED_ST;
      when RX_STARTED_ST =>
                                    if RX_BUSY_HSSL ='0' then -- RX PCS rst is done
                                      rx_pll_pma_started <= '1';
                                    end if;
      when others =>
                                    current_state_rx_pll_pma <= IDLE_ST;
    end case;
  end if;
end process p_rx_pma_pll;

---------------------------------------------------------
-- Process: p_tx_pcs
-- Description: Manages the TX PCS reset of the
--              SpaceFibre HSSL IP
---------------------------------------------------------
p_tx_pcs: process(CLK, RST_N)
begin
  if RST_N ='0' then
    current_state_tx_pcs <= IDLE_ST;
    TX_RST_N_PLIH       <= '0';
    tx_pcs_started       <= '0';
  elsif rising_edge(CLK)  then
    tx_pcs_started       <= '0';
    case current_state_tx_pcs is
      when IDLE_ST =>
                            if pma_pll_seq_end = '1' then -- PMA PLL is locked
                              current_state_tx_pcs <= TX_PULSE_ST;
                            end if;
      when TX_PULSE_ST =>
                            TX_RST_N_PLIH       <= '1'; -- TX PCS rst pulse
                            current_state_tx_pcs <= TX_STARTED_ST;
      when TX_STARTED_ST =>
                            if RX_BUSY_HSSL = '0' then -- TX PCS rst is done
                              tx_pcs_started <= '1';
                            end if;
      when others =>
                            current_state_tx_pcs <= IDLE_ST;
    end case;
  end if;
end process p_tx_pcs;
---------------------------------------------------------
-- Process: p_reset_done
-- Description: Manages HSSL_RESET_DONE_PLIH signal to
--              indicate that the reset of all the IP is done
---------------------------------------------------------
p_reset_done: process(CLK, RST_N)
begin
  if RST_N ='0' then
    HSSL_RESET_DONE_PLIH <= '0';
  elsif rising_edge(CLK)  then
    if tx_pcs_started ='1' and rx_pll_pma_started ='1' then -- TX PCS rst and RX PCS rst are done
      HSSL_RESET_DONE_PLIH <= '1';
    else
      HSSL_RESET_DONE_PLIH <= '0';
    end if;
  end if;
end process p_reset_done;

end architecture rtl;