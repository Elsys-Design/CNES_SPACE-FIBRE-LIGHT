----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2025
--
-- Description : This module describe the Data_word_id_fsm function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library data_link_lib;
use data_link_lib.data_link_lib.all;

entity data_word_id_fsm is
  port (
    RST_N                   : in  std_logic;                                    --! global reset
    CLK                     : in  std_logic;                                    --! Clock generated by GTY IP
		-- data_link_reset (DLRE) interface
    LINK_RESET_DLRE         : in  std_logic;                                    --! Link Reset command
    -- PHY PLUS LANE layer interface
    FIFO_RX_DATA_VALID_PPL  : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    FIFO_RX_RD_EN_DL       : out std_logic;                                   --! Flag to read data in FIFO RX
    DATA_RX_PPL             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    VALID_K_CHARAC_PPL      : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);               --! K charachter valid in the 32-bit DATA_RX_PPL vector
    -- DCCHECK layer interface
    TYPE_FRAME_DWI          : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    NEW_WORD_DWI            : out std_logic;
    END_FRAME_DWI           : out std_logic;
    DATA_DWI                : out std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
		VALID_K_CHARAC_DWI      : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);               --! K charachter valid in the 32-bit DATA_RX_PPL vector
    SEQ_NUM_DWI             : out std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
    CRC_16B_DWI             : out std_logic_vector(15 downto 0);                --! Flag EMPTY of the FIFO RX
    CRC_8B_DWI              : out std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
		MULTIPLIER_DWI          : out std_logic_vector(C_MULT_SIZE-1 downto 0);
		VC_DWI                  : out std_logic_vector(C_CHANNEL_SIZE-1 downto 0);
		RXNOTHING_ACTIVE_DWI    : out std_logic;
    -- OTHER
    CRC_ERR_DCCHECK         : in  std_logic;
    SEQ_ERR_DSCHECK         : in  std_logic;
    FRAME_ERR_DWI           : out std_logic;
		RXERR_DWI               : out std_logic;
		-- MIB
		DATA_COUNTER_RX_DWI     : out  std_logic_vector(6 downto 0);          --! ACK counter RX
		ACK_COUNTER_RX_DWI      : out  std_logic_vector(2 downto 0);          --! ACK counter RX
    NACK_COUNTER_RX_DWI     : out  std_logic_vector(2 downto 0);          --! NACK counter RX
    FCT_COUNTER_RX_DWI      : out  std_logic_vector(3 downto 0);          --! FCT counter RX
    FULL_COUNTER_RX_DWI     : out  std_logic_vector(1 downto 0);          --! FULL counter RX
    RETRY_COUNTER_RX_DWI    : out  std_logic_vector(1 downto 0)           --! RETRY counter RX
  );
end data_word_id_fsm;

architecture rtl of data_word_id_fsm is

----------------------------- Declaration signals -----------------------------

-- Lane Initialisation FSM transition conditions process
   -- Type
type data_word_id_fsm_type is (
   RX_NOTHING_ST,                                                                --! Reset state
   RX_BROADCAST_FRAME_ST,                                                        --! Disabled TX and RX State
   RX_IDLE_FRAME_ST,                                                             --! Waiting State
   RX_DATA_FRAME_ST,                                                             --! Configuration INIT1 State
   RX_BROADCAST_AND_DATA_FRAME_ST
   );
   -- Signals
signal current_state                : data_word_id_fsm_type;                        --! Current state of the Dat Word Identification FSM
signal current_state_r              : data_word_id_fsm_type;                        --! Current state register
signal receiving_frame    : std_logic;
signal type_incom_frame   : std_logic_vector(1 downto 0);
signal data_word_cnt      : unsigned(6 downto 0);
signal bc_word_cnt        : unsigned(1 downto 0);
-- detected signals
signal detected_sdf     : std_logic;
signal detected_edf     : std_logic;
signal detected_sbf     : std_logic;
signal detected_ebf     : std_logic;
signal detected_sif     : std_logic;
signal detected_fct     : std_logic;
signal detected_ack     : std_logic;
signal detected_nack    : std_logic;
signal detected_full    : std_logic;
signal detected_retry   : std_logic;
signal detected_rxerr_i : std_logic;
-- counter signals
signal ack_counter       : unsigned(2 downto 0);
signal nack_counter      : unsigned(2 downto 0);
signal fct_counter       : unsigned(3 downto 0);
signal full_counter      : unsigned(1 downto 0);
signal retry_counter     : unsigned(1 downto 0);

signal toto : std_logic;
begin
	--------------------------------------------------------
	--                  ASSIGNATION
	--------------------------------------------------------
	DATA_COUNTER_RX_DWI  <= std_logic_vector(data_word_cnt);
	ACK_COUNTER_RX_DWI   <= std_logic_vector(ack_counter);
	NACK_COUNTER_RX_DWI  <= std_logic_vector(nack_counter);
	FCT_COUNTER_RX_DWI   <= std_logic_vector(fct_counter);
	FULL_COUNTER_RX_DWI  <= std_logic_vector(full_counter);
	RETRY_COUNTER_RX_DWI <= std_logic_vector(retry_counter);
	RXERR_DWI            <= detected_rxerr_i;
	detected_sdf         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_SDF_WORD   and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- SDF control word detected
	detected_edf         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(7 downto 0)  = C_K28_0_SYMB and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- EDF control word detected
	detected_sbf         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_SBF_WORD   and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- SBF control word detected
	detected_ebf         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(7 downto 0)  = C_K28_2_SYMB and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- EBF control word detected
	detected_sif         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_SIF_WORD   and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- SIF control word detected
	detected_fct         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(7 downto 0)  = C_K28_3_SYMB and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- FCT control word detected
	detected_ack         <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_ACK_WORD   and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- ACK control word detected
	detected_nack        <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_NACK_WORD  and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- NACK control word detected
	detected_full        <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_FULL_WORD  and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- FULL control word detected
	detected_retry       <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL(15 downto 0) = C_RETRY_WORD and VALID_K_CHARAC_PPL = "0001")  else '0';                                   -- RETRY control word detected
	detected_rxerr_i     <= '1' when (FIFO_RX_DATA_VALID_PPL ='1' and DATA_RX_PPL = C_RXERR_WORD              and VALID_K_CHARAC_PPL = "0001" and current_state /= RX_NOTHING_ST) else '0'; -- RXERR control word detected

-------------------------------------------------------------------------------------------
-- Data Word Identification FSM transition conditions process
p_fsm_data_word_id_transition : process(CLK,RST_N)
begin
   if RST_N = '0' then
      current_state          <= RX_NOTHING_ST;
      current_state_r        <= RX_NOTHING_ST;
      FRAME_ERR_DWI          <= '0';
			RXNOTHING_ACTIVE_DWI   <= '0';
   elsif rising_edge(CLK) then
		  FRAME_ERR_DWI         <= '0';
      current_state_r       <= current_state;
			RXNOTHING_ACTIVE_DWI  <= '0';
      case current_state is
         when RX_NOTHING_ST                  => if LINK_RESET_DLRE = '1' then
                                                   current_state  <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                   current_state  <= RX_BROADCAST_FRAME_ST;
                                                elsif detected_sdf ='1' then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_sif ='1' then
                                                   current_state  <= RX_IDLE_FRAME_ST;
                                                end if;
         when RX_DATA_FRAME_ST               => if LINK_RESET_DLRE = '1' or detected_edf = '1' or detected_retry = '1' or CRC_ERR_DCCHECK = '1' or SEQ_ERR_DSCHECK = '1' then
                                                  current_state  <= RX_NOTHING_ST;
				                                        elsif detected_rxerr_i = '1' then
																									RXNOTHING_ACTIVE_DWI   <= '1';
																									current_state         <= RX_NOTHING_ST;
                                                elsif detected_sdf = '1' or detected_sif = '1' or detected_ebf = '1' or data_word_cnt > C_MAX_DATA_FRAME then
																									RXNOTHING_ACTIVE_DWI   <= '1';
                                                  FRAME_ERR_DWI          <= '1';
                                                  current_state          <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                  current_state  <= RX_BROADCAST_AND_DATA_FRAME_ST;
                                                end if;
         when RX_BROADCAST_FRAME_ST          => if LINK_RESET_DLRE = '1' or (detected_ebf = '1' and bc_word_cnt = C_WORD_BC_FRAME) or detected_retry = '1' or CRC_ERR_DCCHECK = '1' or SEQ_ERR_DSCHECK = '1' then
                                                  current_state  <= RX_NOTHING_ST;
				                                        elsif detected_rxerr_i = '1' then
																									RXNOTHING_ACTIVE_DWI  <= '1';
																									current_state         <= RX_NOTHING_ST;
                                                elsif detected_sdf = '1' or detected_sbf = '1' or detected_sif = '1' or detected_edf = '1' or (detected_ebf = '1' and bc_word_cnt /= C_WORD_BC_FRAME) or bc_word_cnt > C_WORD_BC_FRAME then
                                                  RXNOTHING_ACTIVE_DWI  <= '1';
																									FRAME_ERR_DWI         <= '1';
                                                  current_state         <= RX_NOTHING_ST;
                                                end if;

         when RX_BROADCAST_AND_DATA_FRAME_ST => if LINK_RESET_DLRE = '1' or detected_retry = '1' or CRC_ERR_DCCHECK = '1' or SEQ_ERR_DSCHECK = '1' then
                                                  current_state  <= RX_NOTHING_ST;
				                                        elsif detected_rxerr_i = '1' then
																									RXNOTHING_ACTIVE_DWI  <= '1';
																									current_state         <= RX_NOTHING_ST;
                                                elsif (detected_ebf = '1' and bc_word_cnt = C_WORD_BC_FRAME) then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_sdf = '1' or detected_sbf = '1' or detected_sif = '1' or detected_edf = '1' or (detected_ebf = '1' and bc_word_cnt /= C_WORD_BC_FRAME) or bc_word_cnt > C_WORD_BC_FRAME then
                                                  RXNOTHING_ACTIVE_DWI <= '1';
																									FRAME_ERR_DWI        <= '1';
                                                   current_state       <= RX_NOTHING_ST;
                                                end if;

         when RX_IDLE_FRAME_ST               => if LINK_RESET_DLRE = '1' or detected_rxerr_i = '1' or detected_retry = '1' or CRC_ERR_DCCHECK = '1' or SEQ_ERR_DSCHECK = '1' then
                                                  current_state  <= RX_NOTHING_ST;
                                                elsif detected_sbf ='1' then
                                                   current_state  <= RX_BROADCAST_FRAME_ST;
                                                elsif detected_sdf ='1' then
                                                   current_state  <= RX_DATA_FRAME_ST;
                                                elsif detected_edf = '1' or detected_ebf = '1' or data_word_cnt > C_MAX_IDLE_FRAME then
                                                   FRAME_ERR_DWI      <= '1';
                                                   current_state  <= RX_NOTHING_ST;
                                                end if;
         when others                          => current_state  <= RX_NOTHING_ST;
      end case;
   end if;
end process p_fsm_data_word_id_transition;

-- Data Word Identification FSM action on state process
p_comb_state : process(CLK,RST_N)
begin
	if RST_N = '0' then
	  receiving_frame         <= '0';
	  type_incom_frame        <= (others =>'0');
	  data_word_cnt           <= (others =>'0');
	  bc_word_cnt             <= (others =>'0');
	elsif rising_edge(CLK) then
		if current_state = RX_NOTHING_ST then
		  receiving_frame      <= '0';
		  data_word_cnt        <= (others =>'0');
		  bc_word_cnt          <= (others =>'0');
		elsif current_state = RX_DATA_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "01";               -- receiving data frame
		  if (current_state_r = RX_IDLE_FRAME_ST) then
		    data_word_cnt      <= to_unsigned(1,data_word_cnt'length);
		  else
		    data_word_cnt      <= data_word_cnt + 1;
		  end if;
		elsif current_state = RX_BROADCAST_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "10";               -- receiving broadcast frame
		  bc_word_cnt          <= bc_word_cnt + 1;
		  data_word_cnt        <= (others =>'0');
		elsif current_state = RX_BROADCAST_AND_DATA_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "10";               -- receiving broadcast frame
		  bc_word_cnt          <= bc_word_cnt + 1;
		elsif current_state = RX_IDLE_FRAME_ST then
		  receiving_frame      <= '1';
		  type_incom_frame     <= "11";               -- receiving idle frame
		  data_word_cnt        <= data_word_cnt + 1;
		end if;
	end if;
end process p_comb_state;

-- Data Word Identification FSM action on state process
p_data_word_detection : process(CLK,RST_N)
begin
	if RST_N = '0' then
		NEW_WORD_DWI       <= '0';
    SEQ_NUM_DWI        <= (others=> '0');
    CRC_16B_DWI        <= (others=> '0');
    CRC_8B_DWI         <= (others=> '0');
		TYPE_FRAME_DWI     <= (others=> '0');
		DATA_DWI           <= (others=> '0');
		VALID_K_CHARAC_DWI <= (others=> '0');
    END_FRAME_DWI      <= '0';
		MULTIPLIER_DWI     <= (others=> '0');
		VC_DWI             <= (others=> '0');
		ack_counter        <= (others =>'0');
		nack_counter       <= (others =>'0');
		fct_counter        <= (others =>'0');
		full_counter       <= (others =>'0');
		retry_counter      <= (others =>'0');
	elsif rising_edge(CLK) then
    END_FRAME_DWI    <= '0';
		-- Frame treatment
	  if (FIFO_RX_DATA_VALID_PPL ='1') then
			if DATA_RX_PPL(15 downto 0) = C_SDF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SDF control word detected
	  		TYPE_FRAME_DWI     <= C_DATA_FRM;
	  		NEW_WORD_DWI       <= '1';
				DATA_DWI           <= DATA_RX_PPL;
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_0_SYMB and VALID_K_CHARAC_PPL = "0001" and current_state /= RX_NOTHING_ST then -- EDF control word detected
	  		TYPE_FRAME_DWI 		 <= C_DATA_FRM;
	  		NEW_WORD_DWI   		 <= '1';
        END_FRAME_DWI  		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    		 <= DATA_RX_PPL(15 downto 8);
	  		CRC_16B_DWI    		 <= DATA_RX_PPL(31 downto 16);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
	  	elsif DATA_RX_PPL(15 downto 0) = C_SBF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SBF control word detected
	  		TYPE_FRAME_DWI 		 <= C_BC_FRM;
	  		NEW_WORD_DWI   		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_2_SYMB and VALID_K_CHARAC_PPL = "0001" and current_state /= RX_NOTHING_ST then -- EBF control word detected
	  		TYPE_FRAME_DWI		 <= C_BC_FRM;
	  		NEW_WORD_DWI  		 <= '1';
        END_FRAME_DWI 		 <= '1';
				DATA_DWI      		 <= DATA_RX_PPL;
	  		SEQ_NUM_DWI   		 <= DATA_RX_PPL(23 downto 16);
	  		CRC_8B_DWI    		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
	  	elsif DATA_RX_PPL(15 downto 0) = C_SIF_WORD and VALID_K_CHARAC_PPL = "0001" then -- SIF control word detected
	  		TYPE_FRAME_DWI 		 <= C_IDLE_FRM;
	  		NEW_WORD_DWI   		 <= '1';
        END_FRAME_DWI  		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    		 <= DATA_RX_PPL(23 downto 16);
	  		CRC_8B_DWI     		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
	  	elsif DATA_RX_PPL(7 downto 0) = C_K28_3_SYMB and VALID_K_CHARAC_PPL = "0001" then -- FCT control word detected
	  		TYPE_FRAME_DWI 		 <= C_FCT_FRM;
	  		NEW_WORD_DWI   		 <= '1';
        END_FRAME_DWI  		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  		SEQ_NUM_DWI    		 <= DATA_RX_PPL(23 downto 16);
	  		CRC_8B_DWI     		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
				MULTIPLIER_DWI     <= DATA_RX_PPL(15 downto 13);
        VC_DWI             <= DATA_RX_PPL(12 downto 8);
				fct_counter        <= fct_counter + 1;
	  	elsif DATA_RX_PPL(15 downto 0) = C_ACK_WORD and VALID_K_CHARAC_PPL = "0001" then -- ACK control word detected
	  	  TYPE_FRAME_DWI 		 <= C_ACK_FRM;
	  	  NEW_WORD_DWI   		 <= '1';
        END_FRAME_DWI  		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    		 <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
				ack_counter        <= ack_counter + 1;
	  	elsif DATA_RX_PPL(15 downto 0) = C_NACK_WORD and VALID_K_CHARAC_PPL = "0001" then -- NACK control word detected
	  	  TYPE_FRAME_DWI 		 <= C_NACK_FRM;
	  	  NEW_WORD_DWI   		 <= '1';
        END_FRAME_DWI  		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    		 <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
				nack_counter       <= nack_counter + 1;
	  	elsif DATA_RX_PPL(15 downto 0) = C_FULL_WORD and VALID_K_CHARAC_PPL = "0001" then -- FULL control word detected
	  	  TYPE_FRAME_DWI     <= C_FULL_FRM;
	  	  NEW_WORD_DWI       <= '1';
        END_FRAME_DWI      <= '1';
				DATA_DWI           <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI        <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI         <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
				full_counter       <= full_counter + 1;
	  	elsif DATA_RX_PPL(15 downto 0) = C_RETRY_WORD and VALID_K_CHARAC_PPL = "0001" then -- RETRY control word detected
	  	  TYPE_FRAME_DWI 		 <= C_RETRY_FRM;
	  	  NEW_WORD_DWI   		 <= '1';
				DATA_DWI       		 <= DATA_RX_PPL;
	  	  SEQ_NUM_DWI    		 <= DATA_RX_PPL(23 downto 16);
	  	  CRC_8B_DWI     		 <= DATA_RX_PPL(31 downto 24);
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
				retry_counter      <= retry_counter + 1;
	  	elsif DATA_RX_PPL = C_RXERR_WORD and VALID_K_CHARAC_PPL = "0001" then -- RXERR control word detected
        NEW_WORD_DWI   <= '0';
			elsif current_state = RX_IDLE_FRAME_ST or current_state= RX_NOTHING_ST then
					DATA_DWI           <= (others=> '0');
					VALID_K_CHARAC_DWI <= (others=> '0');
					NEW_WORD_DWI       <= '0';
      else
        DATA_DWI           <= DATA_RX_PPL;
				VALID_K_CHARAC_DWI <= VALID_K_CHARAC_PPL;
        NEW_WORD_DWI       <= '1';
	  	end if;
    else
      NEW_WORD_DWI     <= '0';
	  end if;
	end if;
end process p_data_word_detection;

---------------------------------------------------------
-- Process: p_fifo_rd_ppl
-- Description: Write frames into the fifo
---------------------------------------------------------
p_fifo_rd_ppl: process(CLK, RST_N)
begin
	if RST_N = '0' then
		FIFO_RX_RD_EN_DL <= '0';
	elsif rising_edge(CLK) then
		FIFO_RX_RD_EN_DL <= '1';
	end if;
end process p_fifo_rd_ppl;

end architecture rtl;