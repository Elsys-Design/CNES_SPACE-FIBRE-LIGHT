-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 05/08/2025
--
-- Description : This module manages the data writed in the fifo
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_rx_detect_suppr is
  port (
    RST_N                            : in  std_logic;                                          --! global reset
    CLK                              : in  std_logic;                                          --! Clock generated by HSSL IP
    -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
    DATA_RX_PLCWD                    : in std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! 64-bit data from ppl_64_lane_ctrl_word_detect
    VALID_K_CHARAC_PLCWD             : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! 8-bit valid K character flags froml ppl_64_lane_ctrl_word_detect
    DATA_RDY_PLCWD                   : in std_logic_vector(1 downto 0);                        --! Data valid flag ppl_64_lane_ctrl_word_detect
    -- fifo_rx_data (PLFRD) interface
    DATA_RX_PLRDS                    : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! 64-bit data to fifo_rx_data
    VALID_K_CHARAC_PLRDS             : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! 8-bit valid K character flags to fifo_rx_data
    DATA_WR_EN_PLRDS                 : out std_logic                                           --! Data valid flag to fifo_rx_data
  );
end entity;

architecture rtl of ppl_64_rx_detect_suppr is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
type state_type is (
  RX_DATA_1,
  RX_DATA_2
  );

signal current_state       : state_type;

signal data_0              : std_logic_vector(31 downto 0);
signal k_char_0            : std_logic_vector(3 downto 0);

begin

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_detect_suppr
  -- Description: Buffers the data until it has two 32-bit words to write to the fifo
  ---------------------------------------------------------
  p_detect_suppr : process(CLK, RST_N)
  begin
    if RST_N = '0' then
        current_state        <= RX_DATA_1;
        DATA_RX_PLRDS        <= (others => '0');
        VALID_K_CHARAC_PLRDS <= (others => '0');
        DATA_WR_EN_PLRDS     <= '0';
        data_0               <= (others => '0');
        k_char_0             <= (others => '0');
    elsif rising_edge(CLK) then
      case current_state is
          when RX_DATA_1 =>
              if DATA_RDY_PLCWD = "11" then
                DATA_RX_PLRDS        <= DATA_RX_PLCWD;
                VALID_K_CHARAC_PLRDS <= VALID_K_CHARAC_PLCWD;
                DATA_WR_EN_PLRDS     <= '1';
              elsif DATA_RDY_PLCWD = "10" then
                data_0               <= DATA_RX_PLCWD(63 downto 32);
                k_char_0             <= VALID_K_CHARAC_PLCWD(7 downto 4);
                DATA_WR_EN_PLRDS     <= '0';
                current_state        <= RX_DATA_2;
              elsif DATA_RDY_PLCWD = "01" then
                data_0               <= DATA_RX_PLCWD(31 downto 0);
                k_char_0             <= VALID_K_CHARAC_PLCWD(3 downto 0);
                DATA_WR_EN_PLRDS     <= '0';
                current_state        <= RX_DATA_2;
              else
                DATA_WR_EN_PLRDS     <= '0';
              end if;
          when RX_DATA_2 =>
              if DATA_RDY_PLCWD = "11" then
                DATA_RX_PLRDS        <= DATA_RX_PLCWD(31 downto 0) & data_0;
                VALID_K_CHARAC_PLRDS <= VALID_K_CHARAC_PLCWD(3 downto 0) & k_char_0;
                data_0               <= DATA_RX_PLCWD(63 downto 32);
                k_char_0             <= VALID_K_CHARAC_PLCWD(7 downto 4);
                DATA_WR_EN_PLRDS     <= '1';
              elsif DATA_RDY_PLCWD = "10" then
                DATA_RX_PLRDS        <= DATA_RX_PLCWD(63 downto 32) & data_0;
                VALID_K_CHARAC_PLRDS <= VALID_K_CHARAC_PLCWD(7 downto 4) & k_char_0;
                DATA_WR_EN_PLRDS     <= '1';
                current_state        <= RX_DATA_2;
              elsif DATA_RDY_PLCWD = "01" then
                DATA_RX_PLRDS        <= DATA_RX_PLCWD(31 downto 0) & data_0;
                VALID_K_CHARAC_PLRDS <= VALID_K_CHARAC_PLCWD(3 downto 0) & k_char_0;
                DATA_WR_EN_PLRDS     <= '1';
                current_state        <= RX_DATA_2;
              else
                DATA_WR_EN_PLRDS     <= '0';
              end if;
      end case;
    end if;
  end process;
end architecture;

