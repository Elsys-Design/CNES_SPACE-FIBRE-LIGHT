// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_MC_DEFINES_VH
`else
`define B_HBM_MC_DEFINES_VH

// Look-up table parameters
//

`define HBM_MC_ADDR_N  289
`define HBM_MC_ADDR_SZ 32
`define HBM_MC_DATA_SZ 64

// Attribute addresses
//

`define HBM_MC__HBMMC_AP_HINT_MODE    32'h00000000
`define HBM_MC__HBMMC_AP_HINT_MODE_SZ 2

`define HBM_MC__HBMMC_CATTRIP    32'h00000001
`define HBM_MC__HBMMC_CATTRIP_SZ 1

`define HBM_MC__HBMMC_CMD_PAR    32'h00000002
`define HBM_MC__HBMMC_CMD_PAR_SZ 1

`define HBM_MC__HBMMC_CONFIG    32'h00000003
`define HBM_MC__HBMMC_CONFIG_SZ 14

`define HBM_MC__HBMMC_DA28_LOCKOUT    32'h00000004
`define HBM_MC__HBMMC_DA28_LOCKOUT_SZ 1

`define HBM_MC__HBMMC_DATA_ERROR_MODE    32'h00000005
`define HBM_MC__HBMMC_DATA_ERROR_MODE_SZ 3

`define HBM_MC__HBMMC_DQ_RD_PAR    32'h00000006
`define HBM_MC__HBMMC_DQ_RD_PAR_SZ 1

`define HBM_MC__HBMMC_DQ_WR_PAR    32'h00000007
`define HBM_MC__HBMMC_DQ_WR_PAR_SZ 1

`define HBM_MC__HBMMC_DW_LOOPBACK    32'h00000008
`define HBM_MC__HBMMC_DW_LOOPBACK_SZ 1

`define HBM_MC__HBMMC_DW_MISR    32'h00000009
`define HBM_MC__HBMMC_DW_MISR_SZ 3

`define HBM_MC__HBMMC_DW_RD_MUX    32'h0000000a
`define HBM_MC__HBMMC_DW_RD_MUX_SZ 2

`define HBM_MC__HBMMC_ECC    32'h0000000b
`define HBM_MC__HBMMC_ECC_SZ 2

`define HBM_MC__HBMMC_ENTER_SELFREFRESH    32'h0000000c
`define HBM_MC__HBMMC_ENTER_SELFREFRESH_SZ 3

`define HBM_MC__HBMMC_IDLE_TIMEOUT    32'h0000000d
`define HBM_MC__HBMMC_IDLE_TIMEOUT_SZ 27

`define HBM_MC__HBMMC_IDLE_TIMEOUT_EN    32'h0000000e
`define HBM_MC__HBMMC_IDLE_TIMEOUT_EN_SZ 4

`define HBM_MC__HBMMC_INIT_START    32'h0000000f
`define HBM_MC__HBMMC_INIT_START_SZ 20

`define HBM_MC__HBMMC_INT_VREF    32'h00000010
`define HBM_MC__HBMMC_INT_VREF_SZ 3

`define HBM_MC__HBMMC_MAX_PG_IDLE    32'h00000011
`define HBM_MC__HBMMC_MAX_PG_IDLE_SZ 19

`define HBM_MC__HBMMC_MAX_SKIP_CNT    32'h00000012
`define HBM_MC__HBMMC_MAX_SKIP_CNT_SZ 10

`define HBM_MC__HBMMC_MC_DBG_HALT    32'h00000013
`define HBM_MC__HBMMC_MC_DBG_HALT_SZ 3

`define HBM_MC__HBMMC_MC_PM_CAPTURE_TIME    32'h00000014
`define HBM_MC__HBMMC_MC_PM_CAPTURE_TIME_SZ 32

`define HBM_MC__HBMMC_MC_PM_EN    32'h00000015
`define HBM_MC__HBMMC_MC_PM_EN_SZ 16

`define HBM_MC__HBMMC_NA0_BANKADDR_MAP_0    32'h00000016
`define HBM_MC__HBMMC_NA0_BANKADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA0_COLADDR_MAP_0    32'h00000017
`define HBM_MC__HBMMC_NA0_COLADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA0_COLADDR_MAP_1    32'h00000018
`define HBM_MC__HBMMC_NA0_COLADDR_MAP_1_SZ 32

`define HBM_MC__HBMMC_NA0_COLADDR_MAP_2    32'h00000019
`define HBM_MC__HBMMC_NA0_COLADDR_MAP_2_SZ 32

`define HBM_MC__HBMMC_NA0_EXMON_CLR_EXE_CFG_DYN_MCP3    32'h0000001a
`define HBM_MC__HBMMC_NA0_EXMON_CLR_EXE_CFG_DYN_MCP3_SZ 9

`define HBM_MC__HBMMC_NA0_JEDEC_DEVICE_CODE    32'h0000001b
`define HBM_MC__HBMMC_NA0_JEDEC_DEVICE_CODE_SZ 13

`define HBM_MC__HBMMC_NA0_NA_DEST_ID    32'h0000001c
`define HBM_MC__HBMMC_NA0_NA_DEST_ID_SZ 28

`define HBM_MC__HBMMC_NA0_NA_ERR_INJ    32'h0000001d
`define HBM_MC__HBMMC_NA0_NA_ERR_INJ_SZ 32

`define HBM_MC__HBMMC_NA0_NA_NSU_FORCE_ECC_FLIT_ERR    32'h0000001e
`define HBM_MC__HBMMC_NA0_NA_NSU_FORCE_ECC_FLIT_ERR_SZ 32

`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_EN_P0    32'h0000001f
`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_EN_P0_SZ 6

`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_EN_P1    32'h00000020
`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_EN_P1_SZ 6

`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_P0    32'h00000021
`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_P0_SZ 26

`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_P1    32'h00000022
`define HBM_MC__HBMMC_NA0_NA_PM_FILTR_P1_SZ 26

`define HBM_MC__HBMMC_NA0_NA_PM_SMID_FILTR_P0    32'h00000023
`define HBM_MC__HBMMC_NA0_NA_PM_SMID_FILTR_P0_SZ 12

`define HBM_MC__HBMMC_NA0_NA_PM_SMID_FILTR_P1    32'h00000024
`define HBM_MC__HBMMC_NA0_NA_PM_SMID_FILTR_P1_SZ 12

`define HBM_MC__HBMMC_NA0_NA_VC_MAP    32'h00000025
`define HBM_MC__HBMMC_NA0_NA_VC_MAP_SZ 8

`define HBM_MC__HBMMC_NA0_PORT_CONTROL    32'h00000026
`define HBM_MC__HBMMC_NA0_PORT_CONTROL_SZ 26

`define HBM_MC__HBMMC_NA0_RD_CMD_MODE_CFG_MCP    32'h00000027
`define HBM_MC__HBMMC_NA0_RD_CMD_MODE_CFG_MCP_SZ 1

`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_0    32'h00000028
`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_1    32'h00000029
`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_1_SZ 32

`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_2    32'h0000002a
`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_2_SZ 32

`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_3    32'h0000002b
`define HBM_MC__HBMMC_NA0_ROWADDR_MAP_3_SZ 12

`define HBM_MC__HBMMC_NA0_SCRUB_END_ADDRESS    32'h0000002c
`define HBM_MC__HBMMC_NA0_SCRUB_END_ADDRESS_SZ 32

`define HBM_MC__HBMMC_NA0_SCRUB_FREQUENCY    32'h0000002d
`define HBM_MC__HBMMC_NA0_SCRUB_FREQUENCY_SZ 32

`define HBM_MC__HBMMC_NA0_SCRUB_INIT_EN    32'h0000002e
`define HBM_MC__HBMMC_NA0_SCRUB_INIT_EN_SZ 2

`define HBM_MC__HBMMC_NA0_SCRUB_START_ADDRESS    32'h0000002f
`define HBM_MC__HBMMC_NA0_SCRUB_START_ADDRESS_SZ 32

`define HBM_MC__HBMMC_NA0_TGC_CONFIG    32'h00000030
`define HBM_MC__HBMMC_NA0_TGC_CONFIG_SZ 15

`define HBM_MC__HBMMC_NA0_WRCMD_PIPELINE_TIMEOUT_ENABLE_CFG_MCP    32'h00000031
`define HBM_MC__HBMMC_NA0_WRCMD_PIPELINE_TIMEOUT_ENABLE_CFG_MCP_SZ 1

`define HBM_MC__HBMMC_NA0_WRCMD_PIPELINE_TIMEOUT_VALUE_CFG_MCP    32'h00000032
`define HBM_MC__HBMMC_NA0_WRCMD_PIPELINE_TIMEOUT_VALUE_CFG_MCP_SZ 32

`define HBM_MC__HBMMC_NA0_XMPU_CONFIG0_CFG_DYN_MCP3    32'h00000033
`define HBM_MC__HBMMC_NA0_XMPU_CONFIG0_CFG_DYN_MCP3_SZ 5

`define HBM_MC__HBMMC_NA0_XMPU_CONFIG1_CFG_DYN_MCP3    32'h00000034
`define HBM_MC__HBMMC_NA0_XMPU_CONFIG1_CFG_DYN_MCP3_SZ 5

`define HBM_MC__HBMMC_NA0_XMPU_CTRL_CFG_DYN_MCP3    32'h00000035
`define HBM_MC__HBMMC_NA0_XMPU_CTRL_CFG_DYN_MCP3_SZ 4

`define HBM_MC__HBMMC_NA0_XMPU_END_HI0_CFG_DYN_MCP3    32'h00000036
`define HBM_MC__HBMMC_NA0_XMPU_END_HI0_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA0_XMPU_END_HI1_CFG_DYN_MCP3    32'h00000037
`define HBM_MC__HBMMC_NA0_XMPU_END_HI1_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA0_XMPU_END_LO0_CFG_DYN_MCP3    32'h00000038
`define HBM_MC__HBMMC_NA0_XMPU_END_LO0_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA0_XMPU_END_LO1_CFG_DYN_MCP3    32'h00000039
`define HBM_MC__HBMMC_NA0_XMPU_END_LO1_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA0_XMPU_MASTER0_CFG_DYN_MCP3    32'h0000003a
`define HBM_MC__HBMMC_NA0_XMPU_MASTER0_CFG_DYN_MCP3_SZ 26

`define HBM_MC__HBMMC_NA0_XMPU_MASTER1_CFG_DYN_MCP3    32'h0000003b
`define HBM_MC__HBMMC_NA0_XMPU_MASTER1_CFG_DYN_MCP3_SZ 26

`define HBM_MC__HBMMC_NA0_XMPU_START_HI0_CFG_DYN_MCP3    32'h0000003c
`define HBM_MC__HBMMC_NA0_XMPU_START_HI0_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA0_XMPU_START_HI1_CFG_DYN_MCP3    32'h0000003d
`define HBM_MC__HBMMC_NA0_XMPU_START_HI1_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA0_XMPU_START_LO0_CFG_DYN_MCP3    32'h0000003e
`define HBM_MC__HBMMC_NA0_XMPU_START_LO0_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA0_XMPU_START_LO1_CFG_DYN_MCP3    32'h0000003f
`define HBM_MC__HBMMC_NA0_XMPU_START_LO1_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA1_BANKADDR_MAP_0    32'h00000040
`define HBM_MC__HBMMC_NA1_BANKADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA1_COLADDR_MAP_0    32'h00000041
`define HBM_MC__HBMMC_NA1_COLADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA1_COLADDR_MAP_1    32'h00000042
`define HBM_MC__HBMMC_NA1_COLADDR_MAP_1_SZ 32

`define HBM_MC__HBMMC_NA1_COLADDR_MAP_2    32'h00000043
`define HBM_MC__HBMMC_NA1_COLADDR_MAP_2_SZ 32

`define HBM_MC__HBMMC_NA1_EXMON_CLR_EXE_CFG_DYN_MCP3    32'h00000044
`define HBM_MC__HBMMC_NA1_EXMON_CLR_EXE_CFG_DYN_MCP3_SZ 9

`define HBM_MC__HBMMC_NA1_JEDEC_DEVICE_CODE    32'h00000045
`define HBM_MC__HBMMC_NA1_JEDEC_DEVICE_CODE_SZ 13

`define HBM_MC__HBMMC_NA1_NA_DEST_ID    32'h00000046
`define HBM_MC__HBMMC_NA1_NA_DEST_ID_SZ 28

`define HBM_MC__HBMMC_NA1_NA_ERR_INJ    32'h00000047
`define HBM_MC__HBMMC_NA1_NA_ERR_INJ_SZ 32

`define HBM_MC__HBMMC_NA1_NA_NSU_FORCE_ECC_FLIT_ERR    32'h00000048
`define HBM_MC__HBMMC_NA1_NA_NSU_FORCE_ECC_FLIT_ERR_SZ 32

`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_EN_P0    32'h00000049
`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_EN_P0_SZ 6

`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_EN_P1    32'h0000004a
`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_EN_P1_SZ 6

`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_P0    32'h0000004b
`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_P0_SZ 26

`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_P1    32'h0000004c
`define HBM_MC__HBMMC_NA1_NA_PM_FILTR_P1_SZ 26

`define HBM_MC__HBMMC_NA1_NA_PM_SMID_FILTR_P0    32'h0000004d
`define HBM_MC__HBMMC_NA1_NA_PM_SMID_FILTR_P0_SZ 12

`define HBM_MC__HBMMC_NA1_NA_PM_SMID_FILTR_P1    32'h0000004e
`define HBM_MC__HBMMC_NA1_NA_PM_SMID_FILTR_P1_SZ 12

`define HBM_MC__HBMMC_NA1_NA_VC_MAP    32'h0000004f
`define HBM_MC__HBMMC_NA1_NA_VC_MAP_SZ 8

`define HBM_MC__HBMMC_NA1_PORT_CONTROL    32'h00000050
`define HBM_MC__HBMMC_NA1_PORT_CONTROL_SZ 26

`define HBM_MC__HBMMC_NA1_RD_CMD_MODE_CFG_MCP    32'h00000051
`define HBM_MC__HBMMC_NA1_RD_CMD_MODE_CFG_MCP_SZ 1

`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_0    32'h00000052
`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_0_SZ 32

`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_1    32'h00000053
`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_1_SZ 32

`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_2    32'h00000054
`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_2_SZ 32

`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_3    32'h00000055
`define HBM_MC__HBMMC_NA1_ROWADDR_MAP_3_SZ 12

`define HBM_MC__HBMMC_NA1_SCRUB_END_ADDRESS    32'h00000056
`define HBM_MC__HBMMC_NA1_SCRUB_END_ADDRESS_SZ 32

`define HBM_MC__HBMMC_NA1_SCRUB_FREQUENCY    32'h00000057
`define HBM_MC__HBMMC_NA1_SCRUB_FREQUENCY_SZ 32

`define HBM_MC__HBMMC_NA1_SCRUB_INIT_EN    32'h00000058
`define HBM_MC__HBMMC_NA1_SCRUB_INIT_EN_SZ 2

`define HBM_MC__HBMMC_NA1_SCRUB_START_ADDRESS    32'h00000059
`define HBM_MC__HBMMC_NA1_SCRUB_START_ADDRESS_SZ 32

`define HBM_MC__HBMMC_NA1_TGC_CONFIG    32'h0000005a
`define HBM_MC__HBMMC_NA1_TGC_CONFIG_SZ 15

`define HBM_MC__HBMMC_NA1_WRCMD_PIPELINE_TIMEOUT_ENABLE_CFG_MCP    32'h0000005b
`define HBM_MC__HBMMC_NA1_WRCMD_PIPELINE_TIMEOUT_ENABLE_CFG_MCP_SZ 1

`define HBM_MC__HBMMC_NA1_WRCMD_PIPELINE_TIMEOUT_VALUE_CFG_MCP    32'h0000005c
`define HBM_MC__HBMMC_NA1_WRCMD_PIPELINE_TIMEOUT_VALUE_CFG_MCP_SZ 32

`define HBM_MC__HBMMC_NA1_XMPU_CONFIG0_CFG_DYN_MCP3    32'h0000005d
`define HBM_MC__HBMMC_NA1_XMPU_CONFIG0_CFG_DYN_MCP3_SZ 5

`define HBM_MC__HBMMC_NA1_XMPU_CONFIG1_CFG_DYN_MCP3    32'h0000005e
`define HBM_MC__HBMMC_NA1_XMPU_CONFIG1_CFG_DYN_MCP3_SZ 5

`define HBM_MC__HBMMC_NA1_XMPU_CTRL_CFG_DYN_MCP3    32'h0000005f
`define HBM_MC__HBMMC_NA1_XMPU_CTRL_CFG_DYN_MCP3_SZ 4

`define HBM_MC__HBMMC_NA1_XMPU_END_HI0_CFG_DYN_MCP3    32'h00000060
`define HBM_MC__HBMMC_NA1_XMPU_END_HI0_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA1_XMPU_END_HI1_CFG_DYN_MCP3    32'h00000061
`define HBM_MC__HBMMC_NA1_XMPU_END_HI1_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA1_XMPU_END_LO0_CFG_DYN_MCP3    32'h00000062
`define HBM_MC__HBMMC_NA1_XMPU_END_LO0_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA1_XMPU_END_LO1_CFG_DYN_MCP3    32'h00000063
`define HBM_MC__HBMMC_NA1_XMPU_END_LO1_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA1_XMPU_MASTER0_CFG_DYN_MCP3    32'h00000064
`define HBM_MC__HBMMC_NA1_XMPU_MASTER0_CFG_DYN_MCP3_SZ 26

`define HBM_MC__HBMMC_NA1_XMPU_MASTER1_CFG_DYN_MCP3    32'h00000065
`define HBM_MC__HBMMC_NA1_XMPU_MASTER1_CFG_DYN_MCP3_SZ 26

`define HBM_MC__HBMMC_NA1_XMPU_START_HI0_CFG_DYN_MCP3    32'h00000066
`define HBM_MC__HBMMC_NA1_XMPU_START_HI0_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA1_XMPU_START_HI1_CFG_DYN_MCP3    32'h00000067
`define HBM_MC__HBMMC_NA1_XMPU_START_HI1_CFG_DYN_MCP3_SZ 16

`define HBM_MC__HBMMC_NA1_XMPU_START_LO0_CFG_DYN_MCP3    32'h00000068
`define HBM_MC__HBMMC_NA1_XMPU_START_LO0_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NA1_XMPU_START_LO1_CFG_DYN_MCP3    32'h00000069
`define HBM_MC__HBMMC_NA1_XMPU_START_LO1_CFG_DYN_MCP3_SZ 32

`define HBM_MC__HBMMC_NDS    32'h0000006a
`define HBM_MC__HBMMC_NDS_SZ 3

`define HBM_MC__HBMMC_PL    32'h0000006b
`define HBM_MC__HBMMC_PL_SZ 2

`define HBM_MC__HBMMC_RCD_RD    32'h0000006c
`define HBM_MC__HBMMC_RCD_RD_SZ 6

`define HBM_MC__HBMMC_RCD_WR    32'h0000006d
`define HBM_MC__HBMMC_RCD_WR_SZ 6

`define HBM_MC__HBMMC_RD_DBI    32'h0000006e
`define HBM_MC__HBMMC_RD_DBI_SZ 1

`define HBM_MC__HBMMC_REFRESH_MODE    32'h0000006f
`define HBM_MC__HBMMC_REFRESH_MODE_SZ 3

`define HBM_MC__HBMMC_SCAN_VIA_BLI    32'h00000070
`define HBM_MC__HBMMC_SCAN_VIA_BLI_SZ 1

`define HBM_MC__HBMMC_TCCDR    32'h00000071
`define HBM_MC__HBMMC_TCCDR_SZ 6

`define HBM_MC__HBMMC_TCCD_L    32'h00000072
`define HBM_MC__HBMMC_TCCD_L_SZ 6

`define HBM_MC__HBMMC_TCCD_S    32'h00000073
`define HBM_MC__HBMMC_TCCD_S_SZ 6

`define HBM_MC__HBMMC_TCKESR    32'h00000074
`define HBM_MC__HBMMC_TCKESR_SZ 10

`define HBM_MC__HBMMC_TCSR    32'h00000075
`define HBM_MC__HBMMC_TCSR_SZ 1

`define HBM_MC__HBMMC_TEST_MODE    32'h00000076
`define HBM_MC__HBMMC_TEST_MODE_SZ 1

`define HBM_MC__HBMMC_TFAW_L    32'h00000077
`define HBM_MC__HBMMC_TFAW_L_SZ 6

`define HBM_MC__HBMMC_TFAW_S    32'h00000078
`define HBM_MC__HBMMC_TFAW_S_SZ 6

`define HBM_MC__HBMMC_TINIT5    32'h00000079
`define HBM_MC__HBMMC_TINIT5_SZ 10

`define HBM_MC__HBMMC_TMOD    32'h0000007a
`define HBM_MC__HBMMC_TMOD_SZ 10

`define HBM_MC__HBMMC_TMRD    32'h0000007b
`define HBM_MC__HBMMC_TMRD_SZ 10

`define HBM_MC__HBMMC_TRAS    32'h0000007c
`define HBM_MC__HBMMC_TRAS_SZ 6

`define HBM_MC__HBMMC_TRC    32'h0000007d
`define HBM_MC__HBMMC_TRC_SZ 7

`define HBM_MC__HBMMC_TREFI    32'h0000007e
`define HBM_MC__HBMMC_TREFI_SZ 16

`define HBM_MC__HBMMC_TRFC    32'h0000007f
`define HBM_MC__HBMMC_TRFC_SZ 12

`define HBM_MC__HBMMC_TRFCSB    32'h00000080
`define HBM_MC__HBMMC_TRFCSB_SZ 12

`define HBM_MC__HBMMC_TRL    32'h00000081
`define HBM_MC__HBMMC_TRL_SZ 6

`define HBM_MC__HBMMC_TRP    32'h00000082
`define HBM_MC__HBMMC_TRP_SZ 6

`define HBM_MC__HBMMC_TRR    32'h00000083
`define HBM_MC__HBMMC_TRR_SZ 6

`define HBM_MC__HBMMC_TRRD_L    32'h00000084
`define HBM_MC__HBMMC_TRRD_L_SZ 6

`define HBM_MC__HBMMC_TRRD_S    32'h00000085
`define HBM_MC__HBMMC_TRRD_S_SZ 6

`define HBM_MC__HBMMC_TRREFD    32'h00000086
`define HBM_MC__HBMMC_TRREFD_SZ 6

`define HBM_MC__HBMMC_TRTP    32'h00000087
`define HBM_MC__HBMMC_TRTP_SZ 6

`define HBM_MC__HBMMC_TRTW    32'h00000088
`define HBM_MC__HBMMC_TRTW_SZ 6

`define HBM_MC__HBMMC_TWL    32'h00000089
`define HBM_MC__HBMMC_TWL_SZ 5

`define HBM_MC__HBMMC_TWTR_L    32'h0000008a
`define HBM_MC__HBMMC_TWTR_L_SZ 6

`define HBM_MC__HBMMC_TWTR_S    32'h0000008b
`define HBM_MC__HBMMC_TWTR_S_SZ 6

`define HBM_MC__HBMMC_TXP_XS    32'h0000008c
`define HBM_MC__HBMMC_TXP_XS_SZ 27

`define HBM_MC__HBMMC_WR    32'h0000008d
`define HBM_MC__HBMMC_WR_SZ 5

`define HBM_MC__HBMMC_WR_DBI    32'h0000008e
`define HBM_MC__HBMMC_WR_DBI_SZ 1

`define HBM_MC__HBMMC_WTP    32'h0000008f
`define HBM_MC__HBMMC_WTP_SZ 6

`define HBM_MC__SIM_MODEL_TYPE    32'h00000090
`define HBM_MC__SIM_MODEL_TYPE_SZ 24

`define HBM_MC__STACK0_CH1_0_PAGE_HIT    32'h00000091
`define HBM_MC__STACK0_CH1_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH1_0_PHY_ACTIVE    32'h00000092
`define HBM_MC__STACK0_CH1_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH1_0_READ_RATE    32'h00000093
`define HBM_MC__STACK0_CH1_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH1_0_WRITE_RATE    32'h00000094
`define HBM_MC__STACK0_CH1_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH1_1_PAGE_HIT    32'h00000095
`define HBM_MC__STACK0_CH1_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH1_1_PHY_ACTIVE    32'h00000096
`define HBM_MC__STACK0_CH1_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH1_1_READ_RATE    32'h00000097
`define HBM_MC__STACK0_CH1_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH1_1_WRITE_RATE    32'h00000098
`define HBM_MC__STACK0_CH1_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH1_DATA_RATE    32'h00000099
`define HBM_MC__STACK0_CH1_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH2_0_PAGE_HIT    32'h0000009a
`define HBM_MC__STACK0_CH2_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH2_0_PHY_ACTIVE    32'h0000009b
`define HBM_MC__STACK0_CH2_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH2_0_READ_RATE    32'h0000009c
`define HBM_MC__STACK0_CH2_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH2_0_WRITE_RATE    32'h0000009d
`define HBM_MC__STACK0_CH2_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH2_1_PAGE_HIT    32'h0000009e
`define HBM_MC__STACK0_CH2_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH2_1_PHY_ACTIVE    32'h0000009f
`define HBM_MC__STACK0_CH2_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH2_1_READ_RATE    32'h000000a0
`define HBM_MC__STACK0_CH2_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH2_1_WRITE_RATE    32'h000000a1
`define HBM_MC__STACK0_CH2_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH2_DATA_RATE    32'h000000a2
`define HBM_MC__STACK0_CH2_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH3_0_PAGE_HIT    32'h000000a3
`define HBM_MC__STACK0_CH3_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH3_0_PHY_ACTIVE    32'h000000a4
`define HBM_MC__STACK0_CH3_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH3_0_READ_RATE    32'h000000a5
`define HBM_MC__STACK0_CH3_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH3_0_WRITE_RATE    32'h000000a6
`define HBM_MC__STACK0_CH3_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH3_1_PAGE_HIT    32'h000000a7
`define HBM_MC__STACK0_CH3_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH3_1_PHY_ACTIVE    32'h000000a8
`define HBM_MC__STACK0_CH3_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH3_1_READ_RATE    32'h000000a9
`define HBM_MC__STACK0_CH3_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH3_1_WRITE_RATE    32'h000000aa
`define HBM_MC__STACK0_CH3_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH3_DATA_RATE    32'h000000ab
`define HBM_MC__STACK0_CH3_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH4_0_PAGE_HIT    32'h000000ac
`define HBM_MC__STACK0_CH4_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH4_0_PHY_ACTIVE    32'h000000ad
`define HBM_MC__STACK0_CH4_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH4_0_READ_RATE    32'h000000ae
`define HBM_MC__STACK0_CH4_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH4_0_WRITE_RATE    32'h000000af
`define HBM_MC__STACK0_CH4_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH4_1_PAGE_HIT    32'h000000b0
`define HBM_MC__STACK0_CH4_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH4_1_PHY_ACTIVE    32'h000000b1
`define HBM_MC__STACK0_CH4_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH4_1_READ_RATE    32'h000000b2
`define HBM_MC__STACK0_CH4_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH4_1_WRITE_RATE    32'h000000b3
`define HBM_MC__STACK0_CH4_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH4_DATA_RATE    32'h000000b4
`define HBM_MC__STACK0_CH4_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH5_0_PAGE_HIT    32'h000000b5
`define HBM_MC__STACK0_CH5_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH5_0_PHY_ACTIVE    32'h000000b6
`define HBM_MC__STACK0_CH5_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH5_0_READ_RATE    32'h000000b7
`define HBM_MC__STACK0_CH5_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH5_0_WRITE_RATE    32'h000000b8
`define HBM_MC__STACK0_CH5_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH5_1_PAGE_HIT    32'h000000b9
`define HBM_MC__STACK0_CH5_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH5_1_PHY_ACTIVE    32'h000000ba
`define HBM_MC__STACK0_CH5_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH5_1_READ_RATE    32'h000000bb
`define HBM_MC__STACK0_CH5_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH5_1_WRITE_RATE    32'h000000bc
`define HBM_MC__STACK0_CH5_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH5_DATA_RATE    32'h000000bd
`define HBM_MC__STACK0_CH5_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH6_0_PAGE_HIT    32'h000000be
`define HBM_MC__STACK0_CH6_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH6_0_PHY_ACTIVE    32'h000000bf
`define HBM_MC__STACK0_CH6_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH6_0_READ_RATE    32'h000000c0
`define HBM_MC__STACK0_CH6_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH6_0_WRITE_RATE    32'h000000c1
`define HBM_MC__STACK0_CH6_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH6_1_PAGE_HIT    32'h000000c2
`define HBM_MC__STACK0_CH6_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH6_1_PHY_ACTIVE    32'h000000c3
`define HBM_MC__STACK0_CH6_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH6_1_READ_RATE    32'h000000c4
`define HBM_MC__STACK0_CH6_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH6_1_WRITE_RATE    32'h000000c5
`define HBM_MC__STACK0_CH6_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH6_DATA_RATE    32'h000000c6
`define HBM_MC__STACK0_CH6_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH7_0_PAGE_HIT    32'h000000c7
`define HBM_MC__STACK0_CH7_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH7_0_PHY_ACTIVE    32'h000000c8
`define HBM_MC__STACK0_CH7_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH7_0_READ_RATE    32'h000000c9
`define HBM_MC__STACK0_CH7_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH7_0_WRITE_RATE    32'h000000ca
`define HBM_MC__STACK0_CH7_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH7_1_PAGE_HIT    32'h000000cb
`define HBM_MC__STACK0_CH7_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH7_1_PHY_ACTIVE    32'h000000cc
`define HBM_MC__STACK0_CH7_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH7_1_READ_RATE    32'h000000cd
`define HBM_MC__STACK0_CH7_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH7_1_WRITE_RATE    32'h000000ce
`define HBM_MC__STACK0_CH7_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH7_DATA_RATE    32'h000000cf
`define HBM_MC__STACK0_CH7_DATA_RATE_SZ 12

`define HBM_MC__STACK0_CH8_0_PAGE_HIT    32'h000000d0
`define HBM_MC__STACK0_CH8_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH8_0_PHY_ACTIVE    32'h000000d1
`define HBM_MC__STACK0_CH8_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH8_0_READ_RATE    32'h000000d2
`define HBM_MC__STACK0_CH8_0_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH8_0_WRITE_RATE    32'h000000d3
`define HBM_MC__STACK0_CH8_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH8_1_PAGE_HIT    32'h000000d4
`define HBM_MC__STACK0_CH8_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK0_CH8_1_PHY_ACTIVE    32'h000000d5
`define HBM_MC__STACK0_CH8_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK0_CH8_1_READ_RATE    32'h000000d6
`define HBM_MC__STACK0_CH8_1_READ_RATE_SZ 7

`define HBM_MC__STACK0_CH8_1_WRITE_RATE    32'h000000d7
`define HBM_MC__STACK0_CH8_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK0_CH8_DATA_RATE    32'h000000d8
`define HBM_MC__STACK0_CH8_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH1_0_PAGE_HIT    32'h000000d9
`define HBM_MC__STACK1_CH1_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH1_0_PHY_ACTIVE    32'h000000da
`define HBM_MC__STACK1_CH1_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH1_0_READ_RATE    32'h000000db
`define HBM_MC__STACK1_CH1_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH1_0_WRITE_RATE    32'h000000dc
`define HBM_MC__STACK1_CH1_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH1_1_PAGE_HIT    32'h000000dd
`define HBM_MC__STACK1_CH1_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH1_1_PHY_ACTIVE    32'h000000de
`define HBM_MC__STACK1_CH1_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH1_1_READ_RATE    32'h000000df
`define HBM_MC__STACK1_CH1_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH1_1_WRITE_RATE    32'h000000e0
`define HBM_MC__STACK1_CH1_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH1_DATA_RATE    32'h000000e1
`define HBM_MC__STACK1_CH1_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH2_0_PAGE_HIT    32'h000000e2
`define HBM_MC__STACK1_CH2_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH2_0_PHY_ACTIVE    32'h000000e3
`define HBM_MC__STACK1_CH2_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH2_0_READ_RATE    32'h000000e4
`define HBM_MC__STACK1_CH2_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH2_0_WRITE_RATE    32'h000000e5
`define HBM_MC__STACK1_CH2_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH2_1_PAGE_HIT    32'h000000e6
`define HBM_MC__STACK1_CH2_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH2_1_PHY_ACTIVE    32'h000000e7
`define HBM_MC__STACK1_CH2_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH2_1_READ_RATE    32'h000000e8
`define HBM_MC__STACK1_CH2_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH2_1_WRITE_RATE    32'h000000e9
`define HBM_MC__STACK1_CH2_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH2_DATA_RATE    32'h000000ea
`define HBM_MC__STACK1_CH2_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH3_0_PAGE_HIT    32'h000000eb
`define HBM_MC__STACK1_CH3_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH3_0_PHY_ACTIVE    32'h000000ec
`define HBM_MC__STACK1_CH3_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH3_0_READ_RATE    32'h000000ed
`define HBM_MC__STACK1_CH3_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH3_0_WRITE_RATE    32'h000000ee
`define HBM_MC__STACK1_CH3_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH3_1_PAGE_HIT    32'h000000ef
`define HBM_MC__STACK1_CH3_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH3_1_PHY_ACTIVE    32'h000000f0
`define HBM_MC__STACK1_CH3_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH3_1_READ_RATE    32'h000000f1
`define HBM_MC__STACK1_CH3_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH3_1_WRITE_RATE    32'h000000f2
`define HBM_MC__STACK1_CH3_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH3_DATA_RATE    32'h000000f3
`define HBM_MC__STACK1_CH3_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH4_0_PAGE_HIT    32'h000000f4
`define HBM_MC__STACK1_CH4_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH4_0_PHY_ACTIVE    32'h000000f5
`define HBM_MC__STACK1_CH4_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH4_0_READ_RATE    32'h000000f6
`define HBM_MC__STACK1_CH4_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH4_0_WRITE_RATE    32'h000000f7
`define HBM_MC__STACK1_CH4_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH4_1_PAGE_HIT    32'h000000f8
`define HBM_MC__STACK1_CH4_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH4_1_PHY_ACTIVE    32'h000000f9
`define HBM_MC__STACK1_CH4_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH4_1_READ_RATE    32'h000000fa
`define HBM_MC__STACK1_CH4_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH4_1_WRITE_RATE    32'h000000fb
`define HBM_MC__STACK1_CH4_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH4_DATA_RATE    32'h000000fc
`define HBM_MC__STACK1_CH4_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH5_0_PAGE_HIT    32'h000000fd
`define HBM_MC__STACK1_CH5_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH5_0_PHY_ACTIVE    32'h000000fe
`define HBM_MC__STACK1_CH5_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH5_0_READ_RATE    32'h000000ff
`define HBM_MC__STACK1_CH5_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH5_0_WRITE_RATE    32'h00000100
`define HBM_MC__STACK1_CH5_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH5_1_PAGE_HIT    32'h00000101
`define HBM_MC__STACK1_CH5_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH5_1_PHY_ACTIVE    32'h00000102
`define HBM_MC__STACK1_CH5_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH5_1_READ_RATE    32'h00000103
`define HBM_MC__STACK1_CH5_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH5_1_WRITE_RATE    32'h00000104
`define HBM_MC__STACK1_CH5_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH5_DATA_RATE    32'h00000105
`define HBM_MC__STACK1_CH5_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH6_0_PAGE_HIT    32'h00000106
`define HBM_MC__STACK1_CH6_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH6_0_PHY_ACTIVE    32'h00000107
`define HBM_MC__STACK1_CH6_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH6_0_READ_RATE    32'h00000108
`define HBM_MC__STACK1_CH6_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH6_0_WRITE_RATE    32'h00000109
`define HBM_MC__STACK1_CH6_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH6_1_PAGE_HIT    32'h0000010a
`define HBM_MC__STACK1_CH6_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH6_1_PHY_ACTIVE    32'h0000010b
`define HBM_MC__STACK1_CH6_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH6_1_READ_RATE    32'h0000010c
`define HBM_MC__STACK1_CH6_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH6_1_WRITE_RATE    32'h0000010d
`define HBM_MC__STACK1_CH6_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH6_DATA_RATE    32'h0000010e
`define HBM_MC__STACK1_CH6_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH7_0_PAGE_HIT    32'h0000010f
`define HBM_MC__STACK1_CH7_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH7_0_PHY_ACTIVE    32'h00000110
`define HBM_MC__STACK1_CH7_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH7_0_READ_RATE    32'h00000111
`define HBM_MC__STACK1_CH7_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH7_0_WRITE_RATE    32'h00000112
`define HBM_MC__STACK1_CH7_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH7_1_PAGE_HIT    32'h00000113
`define HBM_MC__STACK1_CH7_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH7_1_PHY_ACTIVE    32'h00000114
`define HBM_MC__STACK1_CH7_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH7_1_READ_RATE    32'h00000115
`define HBM_MC__STACK1_CH7_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH7_1_WRITE_RATE    32'h00000116
`define HBM_MC__STACK1_CH7_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH7_DATA_RATE    32'h00000117
`define HBM_MC__STACK1_CH7_DATA_RATE_SZ 12

`define HBM_MC__STACK1_CH8_0_PAGE_HIT    32'h00000118
`define HBM_MC__STACK1_CH8_0_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH8_0_PHY_ACTIVE    32'h00000119
`define HBM_MC__STACK1_CH8_0_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH8_0_READ_RATE    32'h0000011a
`define HBM_MC__STACK1_CH8_0_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH8_0_WRITE_RATE    32'h0000011b
`define HBM_MC__STACK1_CH8_0_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH8_1_PAGE_HIT    32'h0000011c
`define HBM_MC__STACK1_CH8_1_PAGE_HIT_SZ 7

`define HBM_MC__STACK1_CH8_1_PHY_ACTIVE    32'h0000011d
`define HBM_MC__STACK1_CH8_1_PHY_ACTIVE_SZ 64

`define HBM_MC__STACK1_CH8_1_READ_RATE    32'h0000011e
`define HBM_MC__STACK1_CH8_1_READ_RATE_SZ 7

`define HBM_MC__STACK1_CH8_1_WRITE_RATE    32'h0000011f
`define HBM_MC__STACK1_CH8_1_WRITE_RATE_SZ 7

`define HBM_MC__STACK1_CH8_DATA_RATE    32'h00000120
`define HBM_MC__STACK1_CH8_DATA_RATE_SZ 12

`endif  // B_HBM_MC_DEFINES_VH