// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_SNGLBLI_INTF_APB_DEFINES_VH
`else
`define B_HBM_SNGLBLI_INTF_APB_DEFINES_VH

// Look-up table parameters
//

`define HBM_SNGLBLI_INTF_APB_ADDR_N  7
`define HBM_SNGLBLI_INTF_APB_ADDR_SZ 32
`define HBM_SNGLBLI_INTF_APB_DATA_SZ 40

// Attribute addresses
//

`define HBM_SNGLBLI_INTF_APB__CLK_SEL    32'h00000000
`define HBM_SNGLBLI_INTF_APB__CLK_SEL_SZ 40

`define HBM_SNGLBLI_INTF_APB__IS_PCLK_INVERTED    32'h00000001
`define HBM_SNGLBLI_INTF_APB__IS_PCLK_INVERTED_SZ 1

`define HBM_SNGLBLI_INTF_APB__IS_PRESET_N_INVERTED    32'h00000002
`define HBM_SNGLBLI_INTF_APB__IS_PRESET_N_INVERTED_SZ 1

`define HBM_SNGLBLI_INTF_APB__MC_ENABLE    32'h00000003
`define HBM_SNGLBLI_INTF_APB__MC_ENABLE_SZ 40

`define HBM_SNGLBLI_INTF_APB__PHY_ENABLE    32'h00000004
`define HBM_SNGLBLI_INTF_APB__PHY_ENABLE_SZ 40

`define HBM_SNGLBLI_INTF_APB__PHY_PCLK_INVERT    32'h00000005
`define HBM_SNGLBLI_INTF_APB__PHY_PCLK_INVERT_SZ 40

`define HBM_SNGLBLI_INTF_APB__SWITCH_ENABLE    32'h00000006
`define HBM_SNGLBLI_INTF_APB__SWITCH_ENABLE_SZ 40

`endif  // B_HBM_SNGLBLI_INTF_APB_DEFINES_VH