----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2024
--
-- Description : This module checks the validity of the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
use work.data_link_lib.all;

entity data_seq_check is
  port (
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- data_crc_check (DCCHECK) interface
    DATA_DCCHECK           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);        --! Data parallel from Lane Layer
		VALID_K_CHARAC_DCCHECK : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); 
    SEQ_NUM_DCCHECK        : in  std_logic_vector(7 downto 0);                      --! Flag EMPTY of the FIFO RX
    END_FRAME_DCCHECK      : in  std_logic;
    TYPE_FRAME_DCCHECK     : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);  --! Flag EMPTY of the FIFO RX
    NEW_WORD_DCCHECK       : in  std_logic; 
		-- data_err_management (DERRM) interface
		NEAR_END_RPF_DERRM     : in  std_logic; 
		SEQ_NUM_ERR_DSCHECK    : out std_logic;
    -- data_mid_buffer (DMBUF) interface
    DATA_DSCHECK           : out std_logic_vector(C_DATA_LENGTH-1 downto 0);    -- Data write bus
		VALID_K_CHARAC_DSCHECK : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); 
    NEW_WORD_DSCHECK       : out std_logic;                                     -- Write command
    END_FRAME_DSCHECK      : out std_logic;
    FIFO_FULL_DMBUF        : in  std_logic 
  );
end data_seq_check;

architecture rtl of data_seq_check is
---------------------------------------------------------
-----                  Declaration signals          -----
---------------------------------------------------------

signal seq_num_cnt    : unsigned(6 downto 0);   --! Data parallel from Lane Layer
signal seq_num_ok     : std_logic;              --! Data parallel from Lane Layer

begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_seq_num
-- Description: Check the SEQ_NUM for each frame 
---------------------------------------------------------
p_seq_num: process(CLK, RST_N)
begin
	if RST_N = '0' then
	  seq_num_cnt    <= (others => '0'); -- Reset seq_num_cnt	on link reset
		seq_num_ok     <= '0';
    SEQ_NUM_ERR_DSCHECK    <= '0';
	elsif rising_edge(CLK) then
	  if (TYPE_FRAME_DCCHECK = C_DATA_FRM  or TYPE_FRAME_DCCHECK = C_BC_FRM or TYPE_FRAME_DCCHECK = C_FCT_FRM) and END_FRAME_DCCHECK = '1' then
			if SEQ_NUM_DCCHECK /= (NEAR_END_RPF_DERRM & std_logic_vector(seq_num_cnt+1)) then
				SEQ_NUM_ERR_DSCHECK <= '1';
				seq_num_ok  <= '0';
			else
				seq_num_cnt <= seq_num_cnt+1;
				SEQ_NUM_ERR_DSCHECK <= '0';
				seq_num_ok  <= '1';
      end if;
	  elsif (TYPE_FRAME_DCCHECK = C_IDLE_FRM  or TYPE_FRAME_DCCHECK = C_FULL_FRM) and END_FRAME_DCCHECK = '1'then
			if SEQ_NUM_DCCHECK /= (NEAR_END_RPF_DERRM & std_logic_vector(seq_num_cnt)) then
				SEQ_NUM_ERR_DSCHECK <= '1';
				seq_num_ok  <= '0';
			else
				SEQ_NUM_ERR_DSCHECK <= '0';
				seq_num_ok  <= '1';
      end if;
	  end if;
	end if;
end process p_seq_num;
---------------------------------------------------------
-- Process: p_fifo_wr
-- Description: Write frames into the fifo
---------------------------------------------------------
p_fifo_wr: process(CLK, RST_N)
begin
	if RST_N = '0' then
	  DATA_DSCHECK           <= (others => '0');
		VALID_K_CHARAC_DSCHECK <= (others => '0');
		NEW_WORD_DSCHECK       <= '0';
    END_FRAME_DSCHECK      <= '0';
	elsif rising_edge(CLK) then
    END_FRAME_DSCHECK <= END_FRAME_DCCHECK;
		if NEW_WORD_DCCHECK ='1' and FIFO_FULL_DMBUF = '0' then
			NEW_WORD_DSCHECK       <= '1';
			DATA_DSCHECK           <= DATA_DCCHECK;
			VALID_K_CHARAC_DSCHECK <= VALID_K_CHARAC_DCCHECK;
		else
			DATA_DSCHECK           <= (others => '0');
			VALID_K_CHARAC_DSCHECK <= (others => '0');
			NEW_WORD_DSCHECK       <= '0';
		end if;
	end if;
end process p_fifo_wr;

end architecture rtl;