// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_ONE_STACK_INTF_DEFINES_VH
`else
`define B_HBM_ONE_STACK_INTF_DEFINES_VH

// Look-up table parameters
//

`define HBM_ONE_STACK_INTF_ADDR_N  122
`define HBM_ONE_STACK_INTF_ADDR_SZ 32
`define HBM_ONE_STACK_INTF_DATA_SZ 152

// Attribute addresses
//

`define HBM_ONE_STACK_INTF__CLK_SEL_00    32'h00000000
`define HBM_ONE_STACK_INTF__CLK_SEL_00_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_01    32'h00000001
`define HBM_ONE_STACK_INTF__CLK_SEL_01_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_02    32'h00000002
`define HBM_ONE_STACK_INTF__CLK_SEL_02_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_03    32'h00000003
`define HBM_ONE_STACK_INTF__CLK_SEL_03_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_04    32'h00000004
`define HBM_ONE_STACK_INTF__CLK_SEL_04_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_05    32'h00000005
`define HBM_ONE_STACK_INTF__CLK_SEL_05_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_06    32'h00000006
`define HBM_ONE_STACK_INTF__CLK_SEL_06_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_07    32'h00000007
`define HBM_ONE_STACK_INTF__CLK_SEL_07_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_08    32'h00000008
`define HBM_ONE_STACK_INTF__CLK_SEL_08_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_09    32'h00000009
`define HBM_ONE_STACK_INTF__CLK_SEL_09_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_10    32'h0000000a
`define HBM_ONE_STACK_INTF__CLK_SEL_10_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_11    32'h0000000b
`define HBM_ONE_STACK_INTF__CLK_SEL_11_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_12    32'h0000000c
`define HBM_ONE_STACK_INTF__CLK_SEL_12_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_13    32'h0000000d
`define HBM_ONE_STACK_INTF__CLK_SEL_13_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_14    32'h0000000e
`define HBM_ONE_STACK_INTF__CLK_SEL_14_SZ 40

`define HBM_ONE_STACK_INTF__CLK_SEL_15    32'h0000000f
`define HBM_ONE_STACK_INTF__CLK_SEL_15_SZ 40

`define HBM_ONE_STACK_INTF__DATARATE_00    32'h00000010
`define HBM_ONE_STACK_INTF__DATARATE_00_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_01    32'h00000011
`define HBM_ONE_STACK_INTF__DATARATE_01_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_02    32'h00000012
`define HBM_ONE_STACK_INTF__DATARATE_02_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_03    32'h00000013
`define HBM_ONE_STACK_INTF__DATARATE_03_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_04    32'h00000014
`define HBM_ONE_STACK_INTF__DATARATE_04_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_05    32'h00000015
`define HBM_ONE_STACK_INTF__DATARATE_05_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_06    32'h00000016
`define HBM_ONE_STACK_INTF__DATARATE_06_SZ 11

`define HBM_ONE_STACK_INTF__DATARATE_07    32'h00000017
`define HBM_ONE_STACK_INTF__DATARATE_07_SZ 11

`define HBM_ONE_STACK_INTF__DA_LOCKOUT    32'h00000018
`define HBM_ONE_STACK_INTF__DA_LOCKOUT_SZ 40

`define HBM_ONE_STACK_INTF__IS_APB_0_PCLK_INVERTED    32'h00000019
`define HBM_ONE_STACK_INTF__IS_APB_0_PCLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_APB_0_PRESET_N_INVERTED    32'h0000001a
`define HBM_ONE_STACK_INTF__IS_APB_0_PRESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_00_ACLK_INVERTED    32'h0000001b
`define HBM_ONE_STACK_INTF__IS_AXI_00_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_00_ARESET_N_INVERTED    32'h0000001c
`define HBM_ONE_STACK_INTF__IS_AXI_00_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_01_ACLK_INVERTED    32'h0000001d
`define HBM_ONE_STACK_INTF__IS_AXI_01_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_01_ARESET_N_INVERTED    32'h0000001e
`define HBM_ONE_STACK_INTF__IS_AXI_01_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_02_ACLK_INVERTED    32'h0000001f
`define HBM_ONE_STACK_INTF__IS_AXI_02_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_02_ARESET_N_INVERTED    32'h00000020
`define HBM_ONE_STACK_INTF__IS_AXI_02_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_03_ACLK_INVERTED    32'h00000021
`define HBM_ONE_STACK_INTF__IS_AXI_03_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_03_ARESET_N_INVERTED    32'h00000022
`define HBM_ONE_STACK_INTF__IS_AXI_03_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_04_ACLK_INVERTED    32'h00000023
`define HBM_ONE_STACK_INTF__IS_AXI_04_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_04_ARESET_N_INVERTED    32'h00000024
`define HBM_ONE_STACK_INTF__IS_AXI_04_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_05_ACLK_INVERTED    32'h00000025
`define HBM_ONE_STACK_INTF__IS_AXI_05_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_05_ARESET_N_INVERTED    32'h00000026
`define HBM_ONE_STACK_INTF__IS_AXI_05_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_06_ACLK_INVERTED    32'h00000027
`define HBM_ONE_STACK_INTF__IS_AXI_06_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_06_ARESET_N_INVERTED    32'h00000028
`define HBM_ONE_STACK_INTF__IS_AXI_06_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_07_ACLK_INVERTED    32'h00000029
`define HBM_ONE_STACK_INTF__IS_AXI_07_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_07_ARESET_N_INVERTED    32'h0000002a
`define HBM_ONE_STACK_INTF__IS_AXI_07_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_08_ACLK_INVERTED    32'h0000002b
`define HBM_ONE_STACK_INTF__IS_AXI_08_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_08_ARESET_N_INVERTED    32'h0000002c
`define HBM_ONE_STACK_INTF__IS_AXI_08_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_09_ACLK_INVERTED    32'h0000002d
`define HBM_ONE_STACK_INTF__IS_AXI_09_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_09_ARESET_N_INVERTED    32'h0000002e
`define HBM_ONE_STACK_INTF__IS_AXI_09_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_10_ACLK_INVERTED    32'h0000002f
`define HBM_ONE_STACK_INTF__IS_AXI_10_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_10_ARESET_N_INVERTED    32'h00000030
`define HBM_ONE_STACK_INTF__IS_AXI_10_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_11_ACLK_INVERTED    32'h00000031
`define HBM_ONE_STACK_INTF__IS_AXI_11_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_11_ARESET_N_INVERTED    32'h00000032
`define HBM_ONE_STACK_INTF__IS_AXI_11_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_12_ACLK_INVERTED    32'h00000033
`define HBM_ONE_STACK_INTF__IS_AXI_12_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_12_ARESET_N_INVERTED    32'h00000034
`define HBM_ONE_STACK_INTF__IS_AXI_12_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_13_ACLK_INVERTED    32'h00000035
`define HBM_ONE_STACK_INTF__IS_AXI_13_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_13_ARESET_N_INVERTED    32'h00000036
`define HBM_ONE_STACK_INTF__IS_AXI_13_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_14_ACLK_INVERTED    32'h00000037
`define HBM_ONE_STACK_INTF__IS_AXI_14_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_14_ARESET_N_INVERTED    32'h00000038
`define HBM_ONE_STACK_INTF__IS_AXI_14_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_15_ACLK_INVERTED    32'h00000039
`define HBM_ONE_STACK_INTF__IS_AXI_15_ACLK_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__IS_AXI_15_ARESET_N_INVERTED    32'h0000003a
`define HBM_ONE_STACK_INTF__IS_AXI_15_ARESET_N_INVERTED_SZ 1

`define HBM_ONE_STACK_INTF__MC_ENABLE_0    32'h0000003b
`define HBM_ONE_STACK_INTF__MC_ENABLE_0_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_1    32'h0000003c
`define HBM_ONE_STACK_INTF__MC_ENABLE_1_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_2    32'h0000003d
`define HBM_ONE_STACK_INTF__MC_ENABLE_2_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_3    32'h0000003e
`define HBM_ONE_STACK_INTF__MC_ENABLE_3_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_4    32'h0000003f
`define HBM_ONE_STACK_INTF__MC_ENABLE_4_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_5    32'h00000040
`define HBM_ONE_STACK_INTF__MC_ENABLE_5_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_6    32'h00000041
`define HBM_ONE_STACK_INTF__MC_ENABLE_6_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_7    32'h00000042
`define HBM_ONE_STACK_INTF__MC_ENABLE_7_SZ 40

`define HBM_ONE_STACK_INTF__MC_ENABLE_APB    32'h00000043
`define HBM_ONE_STACK_INTF__MC_ENABLE_APB_SZ 40

`define HBM_ONE_STACK_INTF__PAGEHIT_PERCENT_00    32'h00000044
`define HBM_ONE_STACK_INTF__PAGEHIT_PERCENT_00_SZ 7

`define HBM_ONE_STACK_INTF__PHY_ENABLE_00    32'h00000045
`define HBM_ONE_STACK_INTF__PHY_ENABLE_00_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_01    32'h00000046
`define HBM_ONE_STACK_INTF__PHY_ENABLE_01_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_02    32'h00000047
`define HBM_ONE_STACK_INTF__PHY_ENABLE_02_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_03    32'h00000048
`define HBM_ONE_STACK_INTF__PHY_ENABLE_03_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_04    32'h00000049
`define HBM_ONE_STACK_INTF__PHY_ENABLE_04_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_05    32'h0000004a
`define HBM_ONE_STACK_INTF__PHY_ENABLE_05_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_06    32'h0000004b
`define HBM_ONE_STACK_INTF__PHY_ENABLE_06_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_07    32'h0000004c
`define HBM_ONE_STACK_INTF__PHY_ENABLE_07_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_08    32'h0000004d
`define HBM_ONE_STACK_INTF__PHY_ENABLE_08_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_09    32'h0000004e
`define HBM_ONE_STACK_INTF__PHY_ENABLE_09_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_10    32'h0000004f
`define HBM_ONE_STACK_INTF__PHY_ENABLE_10_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_11    32'h00000050
`define HBM_ONE_STACK_INTF__PHY_ENABLE_11_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_12    32'h00000051
`define HBM_ONE_STACK_INTF__PHY_ENABLE_12_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_13    32'h00000052
`define HBM_ONE_STACK_INTF__PHY_ENABLE_13_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_14    32'h00000053
`define HBM_ONE_STACK_INTF__PHY_ENABLE_14_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_15    32'h00000054
`define HBM_ONE_STACK_INTF__PHY_ENABLE_15_SZ 40

`define HBM_ONE_STACK_INTF__PHY_ENABLE_APB    32'h00000055
`define HBM_ONE_STACK_INTF__PHY_ENABLE_APB_SZ 40

`define HBM_ONE_STACK_INTF__PHY_PCLK_INVERT_01    32'h00000056
`define HBM_ONE_STACK_INTF__PHY_PCLK_INVERT_01_SZ 40

`define HBM_ONE_STACK_INTF__READ_PERCENT_00    32'h00000057
`define HBM_ONE_STACK_INTF__READ_PERCENT_00_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_01    32'h00000058
`define HBM_ONE_STACK_INTF__READ_PERCENT_01_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_02    32'h00000059
`define HBM_ONE_STACK_INTF__READ_PERCENT_02_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_03    32'h0000005a
`define HBM_ONE_STACK_INTF__READ_PERCENT_03_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_04    32'h0000005b
`define HBM_ONE_STACK_INTF__READ_PERCENT_04_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_05    32'h0000005c
`define HBM_ONE_STACK_INTF__READ_PERCENT_05_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_06    32'h0000005d
`define HBM_ONE_STACK_INTF__READ_PERCENT_06_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_07    32'h0000005e
`define HBM_ONE_STACK_INTF__READ_PERCENT_07_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_08    32'h0000005f
`define HBM_ONE_STACK_INTF__READ_PERCENT_08_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_09    32'h00000060
`define HBM_ONE_STACK_INTF__READ_PERCENT_09_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_10    32'h00000061
`define HBM_ONE_STACK_INTF__READ_PERCENT_10_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_11    32'h00000062
`define HBM_ONE_STACK_INTF__READ_PERCENT_11_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_12    32'h00000063
`define HBM_ONE_STACK_INTF__READ_PERCENT_12_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_13    32'h00000064
`define HBM_ONE_STACK_INTF__READ_PERCENT_13_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_14    32'h00000065
`define HBM_ONE_STACK_INTF__READ_PERCENT_14_SZ 7

`define HBM_ONE_STACK_INTF__READ_PERCENT_15    32'h00000066
`define HBM_ONE_STACK_INTF__READ_PERCENT_15_SZ 7

`define HBM_ONE_STACK_INTF__SIM_DEVICE    32'h00000067
`define HBM_ONE_STACK_INTF__SIM_DEVICE_SZ 152

`define HBM_ONE_STACK_INTF__STACK_LOCATION    32'h00000068
`define HBM_ONE_STACK_INTF__STACK_LOCATION_SZ 1

`define HBM_ONE_STACK_INTF__SWITCH_ENABLE    32'h00000069
`define HBM_ONE_STACK_INTF__SWITCH_ENABLE_SZ 40

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_00    32'h0000006a
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_00_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_01    32'h0000006b
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_01_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_02    32'h0000006c
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_02_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_03    32'h0000006d
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_03_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_04    32'h0000006e
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_04_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_05    32'h0000006f
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_05_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_06    32'h00000070
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_06_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_07    32'h00000071
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_07_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_08    32'h00000072
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_08_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_09    32'h00000073
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_09_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_10    32'h00000074
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_10_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_11    32'h00000075
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_11_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_12    32'h00000076
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_12_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_13    32'h00000077
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_13_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_14    32'h00000078
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_14_SZ 7

`define HBM_ONE_STACK_INTF__WRITE_PERCENT_15    32'h00000079
`define HBM_ONE_STACK_INTF__WRITE_PERCENT_15_SZ 7

`endif  // B_HBM_ONE_STACK_INTF_DEFINES_VH