-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 05/08/2025
--
-- Description : This module manages the data written in the fifo
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_rx_wr_en_fifo is
  port (
    RST_N                            : in  std_logic;                                   --! Global reset. Active Low
    CLK                              : in  std_logic;                                   --! Clock generated by HSSL IP
    -- ppl_64_lane_ctrl_word_detect (PLCWD) interface
    DATA_RX_PLCWD                    : in std_logic_vector(C_DATA_WIDTH-1 downto 0);    --! 64-bit data from ppl_64_lane_ctrl_word_detect
    VALID_K_CHARAC_PLCWD             : in std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);  --! 8-bit valid K character flags from ppl_64_lane_ctrl_word_detect
    DATA_RDY_PLCWD                   : in std_logic_vector(1 downto 0);                 --! Data valid flag from ppl_64_lane_ctrl_word_detect
    -- fifo_rx_data (PLFRD) interface
    DATA_RX_PLRWEF                    : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to fifo_rx_data
    VALID_K_CHARAC_PLRWEF             : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags to fifo_rx_data
    DATA_RDY_PLRWEF                   : out std_logic_vector(1 downto 0);                --! Data valid flag to fifo_rx_data
    DATA_WR_EN_PLRWEF                 : out std_logic                                    --! Write enable flag to fifo_rx_data
  );
end entity;

architecture rtl of ppl_64_rx_wr_en_fifo is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
begin

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_manage_wr
  --! Manages the data written into the fifo
  ---------------------------------------------------------
  p_manage_wr : process(CLK, RST_N)
  begin
    if RST_N = '0' then
      DATA_RX_PLRWEF        <= (others => '0');
      VALID_K_CHARAC_PLRWEF <= (others => '0');
      DATA_RDY_PLRWEF       <= (others => '0');
      DATA_WR_EN_PLRWEF     <= '0';
    elsif rising_edge(CLK) then
      DATA_RX_PLRWEF        <= DATA_RX_PLCWD;
      VALID_K_CHARAC_PLRWEF <= VALID_K_CHARAC_PLCWD;
      DATA_RDY_PLRWEF       <= DATA_RDY_PLCWD;
      -- At least 1 word is ready
      if DATA_RDY_PLCWD /= "00" then
        DATA_WR_EN_PLRWEF     <= '1';
      -- No word ready
      else
        DATA_WR_EN_PLRWEF     <= '0';
      end if;
    end if;
  end process;
end architecture;

