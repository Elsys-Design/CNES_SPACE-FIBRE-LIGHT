// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSPFP32_DEFINES_VH
`else
`define B_DSPFP32_DEFINES_VH

// Look-up table parameters
//

`define DSPFP32_ADDR_N  31
`define DSPFP32_ADDR_SZ 32
`define DSPFP32_DATA_SZ 64

// Attribute addresses
//

`define DSPFP32__ACASCREG    32'h00000000
`define DSPFP32__ACASCREG_SZ 32

`define DSPFP32__AREG    32'h00000001
`define DSPFP32__AREG_SZ 32

`define DSPFP32__A_FPTYPE    32'h00000002
`define DSPFP32__A_FPTYPE_SZ 24

`define DSPFP32__A_INPUT    32'h00000003
`define DSPFP32__A_INPUT_SZ 56

`define DSPFP32__BCASCSEL    32'h00000004
`define DSPFP32__BCASCSEL_SZ 8

`define DSPFP32__B_D_FPTYPE    32'h00000005
`define DSPFP32__B_D_FPTYPE_SZ 24

`define DSPFP32__B_INPUT    32'h00000006
`define DSPFP32__B_INPUT_SZ 56

`define DSPFP32__FPA_PREG    32'h00000007
`define DSPFP32__FPA_PREG_SZ 32

`define DSPFP32__FPBREG    32'h00000008
`define DSPFP32__FPBREG_SZ 32

`define DSPFP32__FPCREG    32'h00000009
`define DSPFP32__FPCREG_SZ 32

`define DSPFP32__FPDREG    32'h0000000a
`define DSPFP32__FPDREG_SZ 32

`define DSPFP32__FPMPIPEREG    32'h0000000b
`define DSPFP32__FPMPIPEREG_SZ 32

`define DSPFP32__FPM_PREG    32'h0000000c
`define DSPFP32__FPM_PREG_SZ 32

`define DSPFP32__FPOPMREG    32'h0000000d
`define DSPFP32__FPOPMREG_SZ 32

`define DSPFP32__INMODEREG    32'h0000000e
`define DSPFP32__INMODEREG_SZ 32

`define DSPFP32__IS_ASYNC_RST_INVERTED    32'h0000000f
`define DSPFP32__IS_ASYNC_RST_INVERTED_SZ 1

`define DSPFP32__IS_CLK_INVERTED    32'h00000010
`define DSPFP32__IS_CLK_INVERTED_SZ 1

`define DSPFP32__IS_FPINMODE_INVERTED    32'h00000011
`define DSPFP32__IS_FPINMODE_INVERTED_SZ 1

`define DSPFP32__IS_FPOPMODE_INVERTED    32'h00000012
`define DSPFP32__IS_FPOPMODE_INVERTED_SZ 7

`define DSPFP32__IS_RSTA_INVERTED    32'h00000013
`define DSPFP32__IS_RSTA_INVERTED_SZ 1

`define DSPFP32__IS_RSTB_INVERTED    32'h00000014
`define DSPFP32__IS_RSTB_INVERTED_SZ 1

`define DSPFP32__IS_RSTC_INVERTED    32'h00000015
`define DSPFP32__IS_RSTC_INVERTED_SZ 1

`define DSPFP32__IS_RSTD_INVERTED    32'h00000016
`define DSPFP32__IS_RSTD_INVERTED_SZ 1

`define DSPFP32__IS_RSTFPA_INVERTED    32'h00000017
`define DSPFP32__IS_RSTFPA_INVERTED_SZ 1

`define DSPFP32__IS_RSTFPINMODE_INVERTED    32'h00000018
`define DSPFP32__IS_RSTFPINMODE_INVERTED_SZ 1

`define DSPFP32__IS_RSTFPMPIPE_INVERTED    32'h00000019
`define DSPFP32__IS_RSTFPMPIPE_INVERTED_SZ 1

`define DSPFP32__IS_RSTFPM_INVERTED    32'h0000001a
`define DSPFP32__IS_RSTFPM_INVERTED_SZ 1

`define DSPFP32__IS_RSTFPOPMODE_INVERTED    32'h0000001b
`define DSPFP32__IS_RSTFPOPMODE_INVERTED_SZ 1

`define DSPFP32__PCOUTSEL    32'h0000001c
`define DSPFP32__PCOUTSEL_SZ 24

`define DSPFP32__RESET_MODE    32'h0000001d
`define DSPFP32__RESET_MODE_SZ 40

`define DSPFP32__USE_MULT    32'h0000001e
`define DSPFP32__USE_MULT_SZ 64

`endif  // B_DSPFP32_DEFINES_VH