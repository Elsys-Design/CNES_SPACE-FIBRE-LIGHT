`include "B_RFDAC_defines.vh"

reg [`RFDAC_DATA_SZ-1:0] ATTR [0:`RFDAC_ADDR_N-1];
reg [`RFDAC__OPT_CLK_DIST_SZ-1:0] OPT_CLK_DIST_REG = OPT_CLK_DIST;
reg [`RFDAC__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`RFDAC__XPA_ACTIVE_DUTYCYCLE_SZ-1:0] XPA_ACTIVE_DUTYCYCLE_REG = XPA_ACTIVE_DUTYCYCLE;
reg [`RFDAC__XPA_CFG0_SZ-1:0] XPA_CFG0_REG = XPA_CFG0;
reg [`RFDAC__XPA_CFG1_SZ-1:0] XPA_CFG1_REG = XPA_CFG1;
reg [`RFDAC__XPA_CFG2_SZ-1:0] XPA_CFG2_REG = XPA_CFG2;
reg [`RFDAC__XPA_NUM_DACS_SZ-1:0] XPA_NUM_DACS_REG = XPA_NUM_DACS;
reg [`RFDAC__XPA_NUM_DUCS_SZ-1:0] XPA_NUM_DUCS_REG = XPA_NUM_DUCS;
reg [`RFDAC__XPA_PLL_USED_SZ:1] XPA_PLL_USED_REG = XPA_PLL_USED;
reg [`RFDAC__XPA_SAMPLE_RATE_MSPS_SZ-1:0] XPA_SAMPLE_RATE_MSPS_REG = XPA_SAMPLE_RATE_MSPS;

initial begin
  ATTR[`RFDAC__OPT_CLK_DIST] = OPT_CLK_DIST;
  ATTR[`RFDAC__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`RFDAC__XPA_ACTIVE_DUTYCYCLE] = XPA_ACTIVE_DUTYCYCLE;
  ATTR[`RFDAC__XPA_CFG0] = XPA_CFG0;
  ATTR[`RFDAC__XPA_CFG1] = XPA_CFG1;
  ATTR[`RFDAC__XPA_CFG2] = XPA_CFG2;
  ATTR[`RFDAC__XPA_NUM_DACS] = XPA_NUM_DACS;
  ATTR[`RFDAC__XPA_NUM_DUCS] = XPA_NUM_DUCS;
  ATTR[`RFDAC__XPA_PLL_USED] = XPA_PLL_USED;
  ATTR[`RFDAC__XPA_SAMPLE_RATE_MSPS] = XPA_SAMPLE_RATE_MSPS;
end

always @(trig_attr) begin
  OPT_CLK_DIST_REG = ATTR[`RFDAC__OPT_CLK_DIST];
  SIM_DEVICE_REG = ATTR[`RFDAC__SIM_DEVICE];
  XPA_ACTIVE_DUTYCYCLE_REG = ATTR[`RFDAC__XPA_ACTIVE_DUTYCYCLE];
  XPA_CFG0_REG = ATTR[`RFDAC__XPA_CFG0];
  XPA_CFG1_REG = ATTR[`RFDAC__XPA_CFG1];
  XPA_CFG2_REG = ATTR[`RFDAC__XPA_CFG2];
  XPA_NUM_DACS_REG = ATTR[`RFDAC__XPA_NUM_DACS];
  XPA_NUM_DUCS_REG = ATTR[`RFDAC__XPA_NUM_DUCS];
  XPA_PLL_USED_REG = ATTR[`RFDAC__XPA_PLL_USED];
  XPA_SAMPLE_RATE_MSPS_REG = ATTR[`RFDAC__XPA_SAMPLE_RATE_MSPS];
end

// procedures to override, read attribute values

task write_attr;
  input  [`RFDAC_ADDR_SZ-1:0] addr;
  input  [`RFDAC_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`RFDAC_DATA_SZ-1:0] read_attr;
  input  [`RFDAC_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
