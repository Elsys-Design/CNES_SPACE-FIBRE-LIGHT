`include "B_DSP_FP_INMUX_defines.vh"

reg [`DSP_FP_INMUX_DATA_SZ-1:0] ATTR [0:`DSP_FP_INMUX_ADDR_N-1];
reg [`DSP_FP_INMUX__AREG_SZ-1:0] AREG_REG = AREG;
reg [`DSP_FP_INMUX__FPA_PREG_SZ-1:0] FPA_PREG_REG = FPA_PREG;
reg [`DSP_FP_INMUX__FPBREG_SZ-1:0] FPBREG_REG = FPBREG;
reg [`DSP_FP_INMUX__FPDREG_SZ-1:0] FPDREG_REG = FPDREG;
reg [`DSP_FP_INMUX__INMODEREG_SZ-1:0] INMODEREG_REG = INMODEREG;
reg IS_FPINMODE_INVERTED_REG = IS_FPINMODE_INVERTED;
reg IS_RSTFPINMODE_INVERTED_REG = IS_RSTFPINMODE_INVERTED;
reg [`DSP_FP_INMUX__LEGACY_SZ:1] LEGACY_REG = LEGACY;
reg [`DSP_FP_INMUX__RESET_MODE_SZ:1] RESET_MODE_REG = RESET_MODE;
reg [`DSP_FP_INMUX__USE_MULT_SZ:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_FP_INMUX__AREG] = AREG;
  ATTR[`DSP_FP_INMUX__FPA_PREG] = FPA_PREG;
  ATTR[`DSP_FP_INMUX__FPBREG] = FPBREG;
  ATTR[`DSP_FP_INMUX__FPDREG] = FPDREG;
  ATTR[`DSP_FP_INMUX__INMODEREG] = INMODEREG;
  ATTR[`DSP_FP_INMUX__IS_FPINMODE_INVERTED] = IS_FPINMODE_INVERTED;
  ATTR[`DSP_FP_INMUX__IS_RSTFPINMODE_INVERTED] = IS_RSTFPINMODE_INVERTED;
  ATTR[`DSP_FP_INMUX__LEGACY] = LEGACY;
  ATTR[`DSP_FP_INMUX__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_FP_INMUX__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  AREG_REG = ATTR[`DSP_FP_INMUX__AREG];
  FPA_PREG_REG = ATTR[`DSP_FP_INMUX__FPA_PREG];
  FPBREG_REG = ATTR[`DSP_FP_INMUX__FPBREG];
  FPDREG_REG = ATTR[`DSP_FP_INMUX__FPDREG];
  INMODEREG_REG = ATTR[`DSP_FP_INMUX__INMODEREG];
  IS_FPINMODE_INVERTED_REG = ATTR[`DSP_FP_INMUX__IS_FPINMODE_INVERTED];
  IS_RSTFPINMODE_INVERTED_REG = ATTR[`DSP_FP_INMUX__IS_RSTFPINMODE_INVERTED];
  LEGACY_REG = ATTR[`DSP_FP_INMUX__LEGACY];
  RESET_MODE_REG = ATTR[`DSP_FP_INMUX__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_FP_INMUX__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FP_INMUX_ADDR_SZ-1:0] addr;
  input  [`DSP_FP_INMUX_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FP_INMUX_DATA_SZ-1:0] read_attr;
  input  [`DSP_FP_INMUX_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
