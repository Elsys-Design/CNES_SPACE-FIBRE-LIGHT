// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DFE_PRACH_DEFINES_VH
`else
`define B_DFE_PRACH_DEFINES_VH

// Look-up table parameters
//

`define DFE_PRACH_ADDR_N  8
`define DFE_PRACH_ADDR_SZ 32
`define DFE_PRACH_DATA_SZ 64

// Attribute addresses
//

`define DFE_PRACH__ACTIVE_DUTYCYCLE    32'h00000000
`define DFE_PRACH__ACTIVE_DUTYCYCLE_SZ 64

`define DFE_PRACH__CLK_FREQ    32'h00000001
`define DFE_PRACH__CLK_FREQ_SZ 64

`define DFE_PRACH__DECIMATION_RATE    32'h00000002
`define DFE_PRACH__DECIMATION_RATE_SZ 64

`define DFE_PRACH__INCOMING_SAMPLE_RATE    32'h00000003
`define DFE_PRACH__INCOMING_SAMPLE_RATE_SZ 64

`define DFE_PRACH__INCOMING_SAMPLE_RATE_STR    32'h00000004
`define DFE_PRACH__INCOMING_SAMPLE_RATE_STR_SZ 40

`define DFE_PRACH__NUM_ACTIVE_ANTENNAS    32'h00000005
`define DFE_PRACH__NUM_ACTIVE_ANTENNAS_SZ 64

`define DFE_PRACH__NUM_ACTIVE_CHANNELS    32'h00000006
`define DFE_PRACH__NUM_ACTIVE_CHANNELS_SZ 64

`define DFE_PRACH__XPA_CFG0    32'h00000007
`define DFE_PRACH__XPA_CFG0_SZ 16

`endif  // B_DFE_PRACH_DEFINES_VH