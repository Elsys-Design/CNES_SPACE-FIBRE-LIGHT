// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_DSP_OUTPUT58_DEFINES_VH
`else
`define B_DSP_OUTPUT58_DEFINES_VH

// Look-up table parameters
//

`define DSP_OUTPUT58_ADDR_N  11
`define DSP_OUTPUT58_ADDR_SZ 32
`define DSP_OUTPUT58_DATA_SZ 120

// Attribute addresses
//

`define DSP_OUTPUT58__ADREG    32'h00000000
`define DSP_OUTPUT58__ADREG_SZ 32

`define DSP_OUTPUT58__AMULTSEL    32'h00000001
`define DSP_OUTPUT58__AMULTSEL_SZ 16

`define DSP_OUTPUT58__AUTORESET_PATDET    32'h00000002
`define DSP_OUTPUT58__AUTORESET_PATDET_SZ 120

`define DSP_OUTPUT58__AUTORESET_PRIORITY    32'h00000003
`define DSP_OUTPUT58__AUTORESET_PRIORITY_SZ 40

`define DSP_OUTPUT58__BMULTSEL    32'h00000004
`define DSP_OUTPUT58__BMULTSEL_SZ 16

`define DSP_OUTPUT58__DSP_MODE    32'h00000005
`define DSP_OUTPUT58__DSP_MODE_SZ 48

`define DSP_OUTPUT58__IS_RSTP_INVERTED    32'h00000006
`define DSP_OUTPUT58__IS_RSTP_INVERTED_SZ 1

`define DSP_OUTPUT58__LEGACY    32'h00000007
`define DSP_OUTPUT58__LEGACY_SZ 40

`define DSP_OUTPUT58__PREG    32'h00000008
`define DSP_OUTPUT58__PREG_SZ 32

`define DSP_OUTPUT58__RESET_MODE    32'h00000009
`define DSP_OUTPUT58__RESET_MODE_SZ 40

`define DSP_OUTPUT58__USE_MULT    32'h0000000a
`define DSP_OUTPUT58__USE_MULT_SZ 64

`endif  // B_DSP_OUTPUT58_DEFINES_VH