----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2025
--
-- Description : This module describes the top of the Data-Link layer
----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library data_link_lib;
use data_link_lib.data_link_lib.all;

entity data_link is
  generic(
    G_VC_NUM               : integer := 8                                    --! Number of virtual channel
    );
  port(
    RST_N                  : in  std_logic;                              --! global reset
    CLK                    : in  std_logic;                              --! Clock generated by GTY IP
    -- Network layer AXI-Stream TX interface
    AXIS_ARSTN_TX_NW       : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_ACLK_TX_NW        : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_TX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_TX_NW       : in  vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_TX_NW       : in  vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_TX_NW       : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_TX_NW      : in  std_logic_vector(G_VC_NUM downto 0);
    -- Network layer RX interface
    AXIS_ARSTN_RX_NW       : in std_logic_vector(G_VC_NUM downto 0);
    AXIS_ACLK_RX_NW        : in std_logic_vector(G_VC_NUM downto 0);
    AXIS_TREADY_RX_NW      : in  std_logic_vector(G_VC_NUM downto 0);
    AXIS_TDATA_RX_DL       : out vc_data_array(G_VC_NUM downto 0);
    AXIS_TUSER_RX_DL       : out vc_k_array(G_VC_NUM downto 0);
    AXIS_TLAST_RX_DL       : out std_logic_vector(G_VC_NUM downto 0);
    AXIS_TVALID_RX_DL      : out std_logic_vector(G_VC_NUM downto 0);
    CURRENT_TIME_SLOT_NW   : in  std_logic_vector(7 downto 0);          --! Current time slot
    -- Lane layer TX interface
    DATA_TX_DL             : out  std_logic_vector(31 downto 00);         --! Data parallel to be send from Data-Link Layer
    CAPABILITY_TX_DL       : out  std_logic_vector(07 downto 00);         --! Capability send on TX link in INIT3 control word
    NEW_DATA_TX_DL         : out  std_logic;                              --! Flag to write data in FIFO TX
    VALID_K_CHARAC_TX_DL   : out  std_logic_vector(03 downto 00);         --! K charachter valid in the 32-bit DATA_TX_DL vector
    FIFO_TX_FULL_PPL       : in   std_logic;                              --! Flag full of the FIFO TX
    -- Lane layer RX interface
    FIFO_RX_RD_EN_DL        : out  std_logic;                              --! Flag to read data in FIFO RX
    DATA_RX_PPL             : in   std_logic_vector(31 downto 00);         --! Data parallel to be received to Data-Link Layer
    FIFO_RX_EMPTY_PPL       : in   std_logic;                              --! Flag EMPTY of the FIFO RX
    FIFO_RX_DATA_VALID_PPL  : in   std_logic;                              --! Flag DATA_VALID of the FIFO RX
    VALID_K_CHARAC_RX_PPL   : in   std_logic_vector(03 downto 00);         --! K charachter valid in the 32-bit DATA_TR_PPL vector
    FAR_END_CAPA_PPL        : in   std_logic_vector(07 downto 00);         --! Capability field receive in INIT3 control word
    LANE_ACTIVE_PPL         : in  std_logic;                               --! Lane Active flag for the DATA Link Layer
    LANE_RESET_DL           : out std_logic;
    -- MIB  parameters interface
    INTERFACE_RESET_MIB     : in std_logic;                                --! Reset the link and all configuration register of the Data Link layer
    LINK_RESET_MIB          : in std_logic;                                --! Reset the link
    NACK_RST_EN_MIB         : in std_logic;                                --! Enable automatic link reset on NACK reception
    NACK_RST_MODE_MIB       : in std_logic;                                --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
    PAUSE_VC_MIB            : in std_logic_vector(G_VC_NUM downto 0);      --! Pause the corresponding virtual channel after the end of current transmission
    CONTINUOUS_VC_MIB       : in std_logic_vector(G_VC_NUM-1 downto 0);    --! Enable the corresponding virtual channel continuous mode
    -- MIB  status interface
    SEQ_NUMBER_TX_DL        : out std_logic_vector(8-1 downto 0);         --! SEQ_NUMBER in transmission
    SEQ_NUMBER_RX_DL        : out std_logic_vector(8-1 downto 0);         --! SEQ_NUMBER in reception
    CREDIT_VC_DL            : out std_logic_vector(G_VC_NUM-1 downto 0);  --! Indicates if each corresponding far-end input buffer has credit
    INPUT_BUF_OVF_VC_DL     : out std_logic_vector(G_VC_NUM-1 downto 0);
    FCT_CREDIT_OVERFLOW_DL  : out std_logic_vector(G_VC_NUM-1 downto 0);  --! Indicates overflow of each corresponding input buffer
    CRC_LONG_ERROR_DL       : out std_logic;                              --! CRC long error
    CRC_SHORT_ERROR_DL      : out std_logic;                              --! CRC short error
    FRAME_ERROR_DL          : out std_logic;                              --! Frame error
    SEQUENCE_ERROR_DL       : out std_logic;                              --! Sequence error
    FAR_END_LINK_RESET_DL   : out std_logic;                              --! Far-end link reset status
    FRAME_FINISHED_DL       : out std_logic_vector(G_VC_NUM downto 0);    --! Indicates that corresponding channel finished emitting a frame
    FRAME_TX_DL             : out std_logic_vector(G_VC_NUM downto 0);    --! Indicates that corresponding channel is emitting a frame
    DATA_COUNTER_TX_DL      : out std_logic_vector(6 downto 0);           --! Indicate the number of data transmitted in last frame emitted
    DATA_COUNTER_RX_DL      : out std_logic_vector(6 downto 0);           --! Indicate the number of data received in last frame received
    ACK_COUNTER_TX_DL       : out  std_logic_vector(2 downto 0);          --! ACK counter TX
    NACK_COUNTER_TX_DL      : out  std_logic_vector(2 downto 0);          --! NACK counter TX
    FCT_COUNTER_TX_DL       : out  std_logic_vector(3 downto 0);          --! FCT counter TX
    ACK_COUNTER_RX_DL       : out  std_logic_vector(2 downto 0);          --! ACK counter RX
    NACK_COUNTER_RX_DL      : out  std_logic_vector(2 downto 0);          --! NACK counter RX
    FCT_COUNTER_RX_DL       : out  std_logic_vector(3 downto 0);          --! FCT counter RX
    FULL_COUNTER_RX_DL      : out  std_logic_vector(1 downto 0);          --! FULL counter RX
    RETRY_COUNTER_RX_DL     : out  std_logic_vector(1 downto 0);          --! RETRY counter RX
    CURRENT_TIME_SLOT_DL    : out  std_logic_vector(7 downto 0);          --! Current time slot
    RESET_PARAM_DL          : out std_logic;                              --! Reset configuration parameters control
    LINK_RST_ASSERTED_DL    : out std_logic;                              --! Link has been reseted
    NACK_SEQ_NUM_DL         : out std_logic_vector(7 downto 0);           --! NACK Seq_num received
    ACK_SEQ_NUM_DL          : out std_logic_vector(7 downto 0);           --! ACK Seq_num received
    DATA_PULSE_RX_DL        : out std_logic;
    ACK_PULSE_RX_DL         : out std_logic;
    NACK_PULSE_RX_DL        : out std_logic;
    FCT_PULSE_RX_DL         : out std_logic;
    FULL_PULSE_RX_DL        : out std_logic;
    RETRY_PULSE_RX_DL       : out std_logic
  );
end data_link;

architecture Behavioral of data_link is
---------------------------------------------------------
-----                  Module declaration           -----
---------------------------------------------------------
  component data_in_bc_buf is
    port (
    RST_N                  : in  std_logic;                                           --! Global reset (Active-low)
    CLK                    : in  std_logic;                                           --! Global Clock
    -- data_link_reset (DLRE) interface
    LINK_RESET_DLRE        : in  std_logic;                                          --! Link Reset command
    -- AXI-Stream interface
    M_AXIS_ARSTN_NW	       : in  std_logic;                                          --! Active-low asynchronous reset for the AXI-Stream interface
    M_AXIS_ACLK_NW	       : in  std_logic;                                          --! Clock signal for the AXI-Stream interface
    M_AXIS_TVALID_DIBUF	   : out std_logic;                                          --! Indicates that TDATA, TUSER, and TLAST are valid
    M_AXIS_TDATA_DIBUF	   : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! AXI-Stream data bus
    M_AXIS_TLAST_DIBUF	   : out std_logic;                                          --! Indicates the end of a data packet
    M_AXIS_TREADY_NW	     : in  std_logic;                                          --! Receiver ready signal (slave is ready to accept data)
    M_AXIS_TUSER_DIBUF     : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! AXI-Stream user-defined sideband signal
    -- data_desencapsulation_bc (DDESBC) interface
    DATA_DDESBC            : in  std_logic_vector(C_DATA_K_WIDTH-1 downto 0);        --! Data parallel (K character + DATA) from data_desencapsulation_bc
    DATA_EN_DDESBC         : in  std_logic                                           --! Data valid flag associated with DDESBC
  );
  end component;
  component data_in_buf is
    port (
      RST_N                  : in  std_logic;                                          --! Global reset (Active-low)
      CLK                    : in  std_logic;                                          --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        : in  std_logic;                                          --! Link Reset command
      LINK_RESET_DIBUF       : out std_logic;                                          --! Link Reset request to data_link_reset
      -- AXI-Stream interface
      M_AXIS_ARSTN_NW       : in   std_logic;                                          --! Active-low asynchronous reset for the AXI-Stream interface
      M_AXIS_ACLK_NW        : in   std_logic;                                          --! Clock signal for the AXI-Stream interface
      M_AXIS_TVALID_DIBUF   : out  std_logic;                                          --! Indicates that TDATA, TUSER, and TLAST are valid
      M_AXIS_TDATA_DIBUF    : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! AXI-Stream data bus
      M_AXIS_TLAST_DIBUF    : out  std_logic;                                          --! Indicates the end of a data packet
      M_AXIS_TREADY_NW      : in   std_logic;                                          --! Receiver ready signal (slave is ready to accept data)
      M_AXIS_TUSER_DIBUF    : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! AXI-Stream user-defined sideband signal
      -- data_desencapsulation (DDES) interface
      DATA_DDES              : in  std_logic_vector(C_DATA_K_WIDTH-1 downto 0);        --! Data parallel (K character + DATA) from data_desencapsulation
      DATA_EN_DDES           : in  std_logic;                                          --! Data valid flag associated with DATA_DDES
      -- data_mac (DMAC) interface
      REQ_FCT_DIBUF          : out std_logic;                                          --! FCT request to data_mac
      REQ_FCT_DONE_DMAC      : in  std_logic;                                          --! FCT request done flag from data_mac
      --MIB interface
      INPUT_BUF_OVF_DIBUF    : out std_logic                                           --! Input buffer oveflow flag
    );
  end component;

  component data_desencapsulation_bc is
    port (
      CLK                      : in  std_logic;                                    --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        : in std_logic;                                       --! Link Reset command
      -- data_mid_buffer_bc (DMBUFBC)interface
      DATA_DMBUFBC             : in  std_logic_vector(C_DATA_K_WIDTH-1 downto 0);  --! Data parallel (K character + DATA) from data_mid_buffer_bc
      DATA_RD_DDESBC           : out std_logic;                                    --! Read command
      DATA_VALID_DMBUFBC       : in  std_logic;                                    --! Data valid flag associated with DATA_DMBUFBC
      -- data_in_bc_buf (DIBUFBC) interface
      DATA_DDESBC              : out  std_logic_vector(C_DATA_K_WIDTH-1 downto 0); --! Data parallel (K character + DATA) to data_in_bc_buf (BRODACST channel)
      DATA_EN_DDESBC           : out  std_logic                                    --! Data valid flag associated with DATA_DDESBC
    );
  end component;

  component data_desencapsulation is
    generic (
      G_VC_NUM       : integer := 8                                             --! Number of virtual channel
    );
    port (
      CLK                    : in  std_logic;                                   --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        : in std_logic;                                    --! Link Reset command
      -- data_mid_buffer (DMBUF)interface
      DATA_DMBUF             : in  std_logic_vector(C_DATA_K_WIDTH-1 downto 0); --! Data parallel (K character + DATA) from data_mid_buffer
      DATA_RD_DDES           : out std_logic;                                   --! Read command
      DATA_VALID_DMBUF       : in  std_logic;                                   --! Data valid flag associated with DATA_DMBUF
      -- data_in_buf (DIBUF) interface
      DATA_DDES              : out  vc_data_k_array(G_VC_NUM-1 downto 0);       --! Data parallel (K character + DATA) to each data_in_buf (1 per VC)
      DATA_EN_DDES           : out  std_logic_vector(G_VC_NUM-1 downto 0)       --! Data valid flag associated with DATA_DDES
  );
  end component;
  component fifo_dc_drop_bad_frame is
    generic (
      G_DWIDTH                : integer := 8;                                 -- Data bus fifo length
      G_AWIDTH                : integer := 8;                                 -- Address bus fifo length
      G_THRESHOLD_HIGH        : integer := 2**8;                              -- high threshold
      G_THRESHOLD_LOW         : integer := 0                                  -- low threshold
    );
    port (
      RST_N                   : in  std_logic;
      -- Writing port
      WR_CLK                  : in  std_logic;                                -- Clock
      WR_DATA                 : in  std_logic_vector(G_DWIDTH-1 downto 0);    -- Data write bus
      WR_DATA_EN              : in  std_logic;                                -- Write command
      -- Frame control port
      FRAME_ERROR             : in std_logic;                                 -- Valid received data
      END_FRAME               : in std_logic;                                 -- End of frame
      ------------------
      -- Reading port
      RD_CLK                  : in  std_logic;                                -- Clock
      RD_DATA                 : out std_logic_vector(G_DWIDTH-1 downto 0);    -- Data read bus
      RD_DATA_EN              : in  std_logic;                                -- Read command
      RD_DATA_VLD             : out std_logic;                                -- Data valid
      -- Command port
      CMD_FLUSH               : in  std_logic;                                -- fifo flush
      STATUS_BUSY_FLUSH       : out std_logic;                                -- fifo is flushing
      -- Status port
      STATUS_THRESHOLD_HIGH   : out std_logic;                                -- threshold high reached flag (sur WR_CLK)
      STATUS_THRESHOLD_LOW    : out std_logic;                                -- threshold low reached flag (sur RD_CLK)
      STATUS_FULL             : out std_logic;                                -- full fifo flag (sur WR_CLK)
      STATUS_EMPTY            : out std_logic;                                -- empty fifo flag (sur RD_CLK)
      STATUS_LEVEL_WR         : out std_logic_vector(G_AWIDTH-1 downto 0);    -- Niveau de remplissage de la FIFO (sur WR_CLK)
      STATUS_LEVEL_RD         : out std_logic_vector(G_AWIDTH-1 downto 0)     -- Niveau de remplissage de la FIFO (sur RD_CLK)
    );
  end component;

  component data_seq_check is
    port (
      CLK                       : in std_logic;                                           --! Global clock
		  -- data_link_reset (DLRE) interface
		  LINK_RESET_DLRE           : in std_logic;                                           --! Link Reset command
      -- data_crc_check (DCCHECK) interface
      DATA_DCCHECK              : in std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel from data_crc_check
		  VALID_K_CHARAC_DCCHECK    : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K character valid in the 32-bit DATA_DCCHECK vector
		  NEW_WORD_DCCHECK          : in std_logic;                                           --! New word Flag associated with DATA_DCCHECK vector
      END_FRAME_DCCHECK         : in std_logic;                                           --! End frame/control word from data_crc_check
      TYPE_FRAME_DCCHECK        : in std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Current frame/control word type from data_crc_check
      SEQ_NUM_DCCHECK           : in std_logic_vector(7 downto 0);                        --! SEQ_NUM from data_crc_check
		  CRC_ERR_DCCHECK           : in std_logic;                                           --! CRC error flag from data_crc_check
		  FRAME_ERR_DCCHECK         : in std_logic;																					  --! Frame error flag from data_crc_check
		  MULTIPLIER_DCCHECK        : in std_logic_vector(C_MULT_SIZE-1 downto 0);            --! Multiplier value of the current FCT word
		  VC_DCCHECK                : in std_logic_vector(C_CHANNEL_SIZE-1 downto 0);         --! Virtual Channel of the current FCT word
		  RXERR_DCCHECK             : in std_logic;                                           --! RXERR flag detection
      RXERR_ALL_DCCHECK         : in std_logic;                                           --! RXERR flag detection during broadcast and data frame status
		  -- data_err_management (DERRM) interface
		  NEAR_END_RPF_DERRM        : in  std_logic;                                          --! Near-End received polarity flag
		  SEQ_NUM_ACK_DSCHECK       : out std_logic_vector(6 downto 0);                       --! SEQ_NUM ACK value
		  END_FRAME_DSCHECK         : out std_logic;                                          --! End flag of the current frame/control word
		  TYPE_FRAME_DSCHECK        : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);   --! Current frame/control word type
		  TRANS_POL_FLG_DERRM       : in  std_logic;                                          --! Transmission polarity flag
		  CRC_ERR_DSCHECK           : out std_logic;                                          --! CRC error flag for the current frame/control word
		  FRAME_ERR_DSCHECK         : out std_logic;                                          --! Frame error flag for the current frame/control word
		  SEQ_NUM_ERR_DSCHECK       : out std_logic;                                          --! SEQ_NUM error for the current frame/control word
		  RXERR_DSCHECK             : out std_logic;                                          --! RXERR flag for the current frame/control word
      -- data_mid_buffer (DMBUF) interface
      DATA_DSCHECK              : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_mid_buffer (data frame)
		  VALID_K_CHARAC_DSCHECK    : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K character valid in the 32-bit DATA_DSCHECK vector
      NEW_WORD_DSCHECK          : out std_logic;                                          --! New word flag associated with DATA_DSCHECK vector
      END_FRAME_FIFO_DSCHECK    : out std_logic;                                          --! End data frame flag
		  FRAME_ERR_DATA_DSCHECK    : out std_logic;                                          --! Frame error flag for the current data frame
      SEQ_NUM_ERR_DATA_DSCHECK  : out std_logic;                                          --! SEQ_NUM error for the current data frame
      CRC_ERR_DATA_DSCHECK      : out std_logic;                                          --! CRC error flag for the current data frame
		  RXERR_DATA_DSCHECK        : out std_logic;                                          --! RXERR flag for the current data frame
		  -- data_mid_buffer_bc (DMBUFBC) interface
		  DATA_BC_DSCHECK           : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_mid_buffer_bc (broadcast frame)
		  VALID_K_CHARAC_BC_DSCHECK : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K character valid in the 32-bit DATA_BC_DSCHECK vector
      NEW_WORD_BC_DSCHECK       : out std_logic;                                          --! New word flag associated with DATA_BC_DSCHECK vector
      END_FRAME_FIFO_BC_DSCHECK : out std_logic;                                          --! End broadcast frame flag
		  FRAME_ERR_BC_DSCHECK      : out std_logic;                                          --! Frame error flag for the current broadcast frame
		  SEQ_NUM_ERR_BC_DSCHECK    : out std_logic;                                          --! SEQ_NUM error for the current broadcast frame
		  CRC_ERR_BC_DSCHECK        : out std_logic;                                          --! CRC error flag for the current broadcast frame
		  RXERR_BC_DSCHECK          : out std_logic;                                          --! RXERR flag for the current broadcast frame
		  -- data_out_buff (DOBUF) interface
		  FCT_FAR_END_DSCHECK       : out std_logic_vector(C_VC_NUM-1 downto 0);              --! FCT received flag for each virtual channel
		  M_VAL_DSCHECK             : out std_logic_vector(C_M_SIZE-1 downto 0);              --! M value associated with FCT_FAR_END_DSCHECK
		  -- MIB
		  SEQ_NUM_DSCHECK           : out std_logic_vector(7 downto 0);                       --! last SEQ_NUM
		  NACK_SEQ_NUM_DSCHECK      : out std_logic_vector(7 downto 0);                       --! last NACK SEQ_NUM
      ACK_SEQ_NUM_DSCHECK       : out std_logic_vector(7 downto 0);                       --! last ACK SEQ_NUM
		  ACK_COUNTER_RX_DSCHECK    : out std_logic_vector(2 downto 0);                       --! ACK counter RX
      NACK_COUNTER_RX_DSCHECK   : out std_logic_vector(2 downto 0);                       --! NACK counter RX
      FCT_COUNTER_RX_DSCHECK    : out std_logic_vector(3 downto 0);                       --! FCT counter RX
      FULL_COUNTER_RX_DSCHECK   : out std_logic_vector(1 downto 0);                       --! FULL counter RX
		  ACK_PULSE_RX_DSCHECK      : out std_logic;                                          --! New ACK received flag
		  NACK_PULSE_RX_DSCHECK     : out std_logic;                                          --! New NACK received flag
		  FCT_PULSE_RX_DSCHECK      : out std_logic;                                          --! New FCT received flag
		  FULL_PULSE_RX_DSCHECK     : out std_logic                                           --! New FULL received flag
  );
  end component;

  component data_crc_check is
    port (
      CLK                    : in  std_logic;                                           --! Global clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        : in std_logic;                                            --! Link Reset command
      -- data_word_identification (DWI) interface
      DATA_DWI               : in std_logic_vector(C_DATA_LENGTH-1 downto 0);           --! Data parallel from data_word_id_fsm
      VALID_K_CHARAC_DWI     : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);   --! K character valid in the 32-bit DATA_DWI vector
      NEW_WORD_DWI           : in std_logic;                                            --! New word Flag from data_word_id_fsm
      END_FRAME_DWI          : in std_logic;                                            --! End frame/control word from data_word_id_fsm
      SEQ_NUM_DWI            : in std_logic_vector(7 downto 0);                         --! SEQ_NUM from data_word_id_fsm
      CRC_16B_DWI            : in std_logic_vector(15 downto 0);                        --! 16-bit CRC (data frame)  from data_word_id_fsm
      CRC_8B_DWI             : in std_logic_vector(7 downto 0);                         --! 8-bit CRC from data_word_id_fsm
      TYPE_FRAME_DWI         : in std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);     --! Current frame/control word type from data_word_id_fsm
      FRAME_ERR_DWI          : in std_logic;                                            --! Frame error flag from data_word_id_fsm
      MULTIPLIER_DWI         : in std_logic_vector(C_MULT_SIZE-1 downto 0);             --! Multiplier value of the current FCT word
		  VC_DWI                 : in std_logic_vector(C_CHANNEL_SIZE-1 downto 0);          --! Virtual Channel of the current FCT word
      RXERR_DWI              : in std_logic;                                            --! RXERR flag detection
		  RXERR_ALL_DWI          : in std_logic;                                            --! RXERR flag detection during broadcast and data frame status
      RXNOTHING_ACTIVE_DWI   : in std_logic;                                            --! RXNOTHING state of the data_word_id_fsm flag
      -- data_seq_check (DSCHECK) interface
      NEW_WORD_DCCHECK       : out std_logic;                                           --! New word flag associated with DATA_DCCHECK
      DATA_DCCHECK           : out std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel to data_seq_check
      VALID_K_CHARAC_DCCHECK : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K character valid in the 32-bit DATA_DCCHECK vector
      END_FRAME_DCCHECK      : out std_logic;                                           --! End frame/control word flag
      TYPE_FRAME_DCCHECK     : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Current frame/control word type
      SEQ_NUM_DCCHECK        : out std_logic_vector(7 downto 0);                        --! SEQ_NUM value
      CRC_ERR_DCCHECK        : out std_logic;                                           --! CRC error flag
      FRAME_ERR_DCCHECK      : out std_logic;                                           --! Frame error flag for the current frame
      MULTIPLIER_DCCHECK     : out std_logic_vector(C_MULT_SIZE-1 downto 0);            --! Multiplier value of the current FCT word
		  VC_DCCHECK             : out std_logic_vector(C_CHANNEL_SIZE-1 downto 0);         --! Virtual Channel of the current FCT word
      RXERR_DCCHECK          : out std_logic;                                           --! RXERR flag for the current frame
      RXERR_ALL_DCCHECK      : out std_logic;                                           --! RXERR flag during broadcast and data frame status
      -- MIB
      CRC_LONG_ERR_DCCHECK   : out std_logic;                                           --! CRC 16-bit error flag
      CRC_SHORT_ERR_DCCHECK  : out std_logic                                            --! CRC 8-bit error flag
  );
  end component;

  component data_word_id_fsm is
    port (
      CLK                     : in  std_logic;                                           --! Global clock
		  -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE         : in  std_logic;                                           --! Link Reset command
      -- PHY PLUS LANE layer interface
      FIFO_RX_DATA_VALID_PPL  : in  std_logic;                                           --! Flag DATA_VALID of the FIFO RX from Lane layer
      FIFO_RX_RD_EN_DL       : out std_logic;                                            --! Flag to read data in FIFO RX
      DATA_RX_PPL             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel from Lane Layer
      VALID_K_CHARAC_PPL      : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K character valid in the 32-bit DATA_RX_PPL vector
      -- data_crc_check (DCCHECK) interface
      TYPE_FRAME_DWI          : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);     --! Current frame/control word type
      NEW_WORD_DWI            : out std_logic;                                            --! New word flag associated to DATA_DWI
      END_FRAME_DWI           : out std_logic;                                            --! End frame/control word flag
      DATA_DWI                : out std_logic_vector(C_DATA_LENGTH-1 downto 0);           --! Data parallel to data_crc_check
		  VALID_K_CHARAC_DWI      : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K character valid in the 32-bit DATA_DWI vector
      SEQ_NUM_DWI             : out std_logic_vector(7 downto 0);                 				--! SEQ_NUM of the current control word
      CRC_16B_DWI             : out std_logic_vector(15 downto 0);                				--! 16-bit CRC (data frame)  of the current control word
      CRC_8B_DWI              : out std_logic_vector(7 downto 0);                 				--! 8-bit CRC of the current control word
		  MULTIPLIER_DWI          : out std_logic_vector(C_MULT_SIZE-1 downto 0);     				--! Multiplier value of the current FCT word
		  VC_DWI                  : out std_logic_vector(C_CHANNEL_SIZE-1 downto 0);  				--! Virtual Channel of the current FCT word
		  RXNOTHING_ACTIVE_DWI    : out std_logic;                                  					--! RXNOTHING state of the data_word_id_fsm flag
		  RXERR_DWI               : out std_logic; 																						--! RXERR flag detection
		  RXERR_ALL_DWI           : out std_logic; 																						--! RXERR flag detection during broadcast and data frame status
      -- Error interface
      CRC_ERR_DCCHECK         : in  std_logic;                                            --! CRC error flag from data_crc_check
      SEQ_ERR_DSCHECK         : in  std_logic;                                            --! SEQ_NUM error flag from data_seq_check
      FRAME_ERR_DWI           : out std_logic;                                            --! Frame error flag
		  -- MIB
		  DATA_COUNTER_RX_DWI     : out  std_logic_vector(6 downto 0);                        --! Data counter RX
      RETRY_COUNTER_RX_DWI    : out  std_logic_vector(1 downto 0);                        --! RETRY counter RX
		  DATA_PULSE_RX_DWI       : out std_logic;                                            --! New data received flag
		  RETRY_PULSE_RX_DWI      : out std_logic                                             --! New RETRY received flag
    );
  end component;

  component data_link_reset is
    generic (
      G_VC_NUM       : integer := 8                                        --! Number of virtual channels
    );
    port (
      RST_N                   : in  std_logic;                              --! Global reset (Active-low)
      CLK                     : in  std_logic;                              --! Global clock
      -- Link Reset
      LINK_RESET_DLRE         : out std_logic;                              --! Link Reset command
      -- data_in_buf (DIBUF) interface
      LINK_RESET_DIBUF        : in  std_logic_vector(G_VC_NUM-1 downto 0);  --! Link Reset request from data_in_buf
      -- data_err_management (DERRM) interface
      LINK_RESET_DERRM        : in std_logic;                               --! Link Reset request from data_err_management
      -- Lane interface
      LANE_RESET_DLRE         : out std_logic;                              --! Lane Reset command
      NEAR_END_CAPA_DLRE      : out std_logic_vector(7 downto 0);           --! Near-end capability
      LANE_ACTIVE_PPL         : in  std_logic;                              --! Lane active flag
      FAR_END_CAPA_PPL        : in  std_logic_vector(7 downto 0);           --! Far-end capability
      --MIB interface
      RESET_PARAM_DLRE        : out std_logic;                              --! Reset all MIB parameters command
      INTERFACE_RESET_MIB     : in  std_logic;                              --! Interface Reset request
      LINK_RESET_MIB          : in  std_logic                               --! Link Reset request
    );
  end component;
  component data_err_management is
    port (
      CLK                      : in std_logic;                                --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE          : in  std_logic;                               --! Link Reset command
      LINK_RESET_DERRM         : out std_logic;                               --! Link Reset request
      -- data_seq_check (DSCHECK) interface
      TYPE_FRAME_DSCHECK       : in std_logic_vector(3 downto 0);             --! Current frame/control word type from data_seq_check
      END_FRAME_DSCHECK        : in std_logic;                                --! End flag of the current frame/control word from data_seq_check
      SEQ_ERR_DSCHECK          : in std_logic;                                --! SEQ_NUM error for the current frame/control word from data_seq_check
      SEQ_NUM_ACK_DSCHECK      : in std_logic_vector(6 downto 0);             --! SEQ_NUM ACK value from data_seq_check
      FAR_END_RPF_DSCHECK      : in std_logic;                                --! Far-end RPF flag
      NEAR_END_RPF_DERRM       : out std_logic;                               --! Near-end RPF flag
      CRC_ERR_DSCHECK          : in std_logic;                                --! CRC error flag for the current frame/control word from data_seq_check
      FRAME_ERR_DSCHECK        : in std_logic;                                --! Frame error flag for the current frame/control word from data_seq_check
      RXERR_DSCHECK            : in std_logic;                                --! Receive error flag from data_word_interface
      -- data_mac (DMAC) interface
      REQ_ACK_DERRM            : out std_logic;                               --! ACK request to data_mac
      REQ_NACK_DERRM           : out std_logic;                               --! NACK request to data_mac
      TRANS_POL_FLG_DERRM      : out std_logic;                               --! Transmission polarity flag to data_mac
      SEQ_NUM_ACK_DERRM        : out std_logic_vector(7 downto 0);            --! SEQ_NUM ACK value to data_mac
      REQ_ACK_DONE_DMAC        : in std_logic;                                --! Acknowledge done signal from data_mac
      -- MIB  interface
      NACK_RST_EN_MIB          : in std_logic;                                --! Enable automatic link reset on NACK reception
      NACK_RST_MODE_MIB        : in std_logic                                 --! Up for instant link reset on NACK reception, down for link reset at the end of the current received frame on NACK reception
  );
    end component;
  component data_out_bc_buf is
    port (
      RST_N                 : in  std_logic;                                          --! Global reset (Active-low)
      CLK                   : in  std_logic;                                          --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        :in  std_logic;                                          --! Link Reset command
      -- AXI-Stream interface
      S_AXIS_ARSTN_NW	      : in std_logic;                                           --! Active-low asynchronous reset for the AXI-Stream interface
		  S_AXIS_ACLK_NW	      : in std_logic;                                           --! Clock signal for the AXI-Stream interface
		  S_AXIS_TREADY_DL      : out std_logic;                                          --! Indicates that TDATA, TUSER, and TLAST are valid
		  S_AXIS_TDATA_NW       : in std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! AXI-Stream data bus
		  S_AXIS_TUSER_NW       : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! Indicates the end of a data packet
		  S_AXIS_TLAST_NW       : in std_logic;                                           --! Receiver ready signal (slave is ready to accept data)
		  S_AXIS_TVALID_NW      : in std_logic;                                           --! AXI-Stream user-defined sideband signal
      -- data_mac (DMAC) interface
      VC_READY_DOBUF        : out  std_logic;                                          --! Virtual Channel ready flag
      DATA_DOBUF            : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_mac
      VALID_K_CHARAC_DOBUF  : out  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K character valid in the 32-bit DATA_DOBUF vector
      DATA_VALID_DOBUF      : out  std_logic;                                          --! Data valid flag associated with DATA_DOBUF
      END_PACKET_DOBUF      : out  std_logic;                                          --! End packet flag
      VC_RD_EN_DMAC         : in   std_logic                                           --! Read command from data_mac
    );
  end component;
  component data_out_buff is
    port (
      RST_N                 : in  std_logic;                                          --! Global reset (Active-low)
      CLK                   : in  std_logic;                                          --! Global Clock
      -- phy_plus_lane (PPL) interface
      LANE_ACTIVE_ST_PPL    : in  std_logic;                                          --! Lane Active state flag
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        :in  std_logic;                                          --! Link Reset command
      -- AXI-Stream interface
      S_AXIS_ARSTN_NW	      : in  std_logic;                                          --! Active-low asynchronous reset signal for the AXI-Stream i
		  S_AXIS_ACLK_NW	      : in  std_logic;                                          --! Clock signal for the AXI-Stream interface
		  S_AXIS_TREADY_DL      : out std_logic;                                          --! Ready signal from the slave indicating it can accept data
		  S_AXIS_TDATA_NW       : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data bus carrying the actual payload
		  S_AXIS_TUSER_NW       : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! User-defined sideband information (optional)
		  S_AXIS_TLAST_NW       : in  std_logic;                                          --! Signal indicating the last transfer in a packet
		  S_AXIS_TVALID_NW      : in  std_logic;                                          --! Valid signal indicating that the data on TDATA is valid
      -- data_mac (DMAC) interface
      VC_READY_DOBUF        : out std_logic;                                          --! Virtual Channel ready flag
      DATA_DOBUF            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_mac
      VALID_K_CHARAC_DOBUF  : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K character valid in the 32-bit DATA_DOBUF vector
      DATA_VALID_DOBUF      : out std_logic;                                          --! Data valid flag associated with DATA_DOBUF
      END_PACKET_DOBUF      : out std_logic;                                          --! End packet flag
      VC_RD_EN_DMAC         : in  std_logic;                                          --! Read command from data_mac
      --DSCHECK interface
      M_VAL_DSCHECK         : in  std_logic_vector(C_M_SIZE-1 downto 0);              --! M value associated with FCT_FAR_END_DSCHECK
      FCT_FAR_END_DSCHECK   : in  std_logic;                                          --! FCT Fare-end received flag
      --MIB Interface
      FCT_CC_OVF_DOBUF      : out std_logic;                                          --! FCT credit counter overflow flag
      CREDIT_VC_DOBUF       : out std_logic;                                          --! Has credit flag (crdit counter > 0)
      VC_CONT_MODE_MIB      : in  std_logic                                           --! Continuous mode command
    );
  end component;

  component data_mac is
    generic(
      G_VC_NUM           : integer := 8                                              --! Number of virtual channel
      );
    port (
      CLK                  : in  std_logic;                                          --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE        :in  std_logic;                                         --! Link Reset command
      -- phy_plus_lane (PPL) interface
      LANE_ACTIVE_PPL      : in  std_logic;                                          --! Lane Active flag for the DATA Link Layer
      -- data_err_management (DERRM) interface
      REQ_ACK_DERRM        : in  std_logic;                                          --! ACK request from data_err_management
      REQ_NACK_DERRM       : in  std_logic;                                          --! NACK request from data_err_management
      TRANS_POL_FLG_DERRM  : in  std_logic;                                          --! Transmission polarity flag from data_err_management
      REQ_ACK_DONE_DMAC    : out std_logic;                                          --! Acknowledge done signal to data_err_management
      SEQ_NUM_ACK_DERRM    : in  std_logic_vector(7 downto 0);                       --! SEQ_NUM ACK value from data_err_management
      -- data_in_buf (DIBUF) interface
      REQ_FCT_DIBUF        : in  std_logic_vector(G_VC_NUM-1 downto 0);              --! FCT request from data_in_buf
      REQ_FCT_DONE_DMAC    : out std_logic_vector(G_VC_NUM-1 downto 0);              --! FCT request done flag to data_in_buf
      -- data_out_buff (DOBUF) interface
      VC_READY_DOBUF       : in  std_logic_vector(G_VC_NUM downto 0);                --! Virtual Channel ready flag vector
      VC_DATA_DOBUF        : in  vc_data_array(G_VC_NUM downto 0);                   --! Array of data vector for each Virtual Channel
      VC_VALID_K_CHAR_DOBUF: in  vc_k_array(G_VC_NUM downto 0);                      --! Array of K character valid in the 32-bit VC_DATA_DOBUF
      VC_DATA_VALID_DOBUF  : in  std_logic_vector(G_VC_NUM downto 0);                --! Data valid flag associated with VC_DATA_DOBUF
      VC_END_PACKET_DOBUF  : in  std_logic_vector(G_VC_NUM downto 0);                --! End packet flag vector for each Virtual Channel
      VC_RD_EN_DMAC        : out  std_logic_vector(G_VC_NUM downto 0);               --! Read command vector for each Virtual Channel
      -- MIB interface
      VC_PAUSE_MIB         : in  std_logic_vector(G_VC_NUM downto 0);                --! Pause the corresponding virtual channel after the end of current transmission
      VC_END_EMISSION_DMAC : out std_logic_vector(G_VC_NUM downto 0);                --! Indicates that corresponding channel finished emitting a frame
      VC_RUN_EMISSION_DMAC : out std_logic_vector(G_VC_NUM downto 0);                --! Indicates that corresponding channel is emitting a frame
      DATA_COUNTER_TX_DMAC : out std_logic_vector(6 downto 0);                       --! Indicate the number of data transmitted in last frame emitted
      ACK_COUNTER_TX_DMAC  : out  std_logic_vector(2 downto 0);                      --! ACK counter TX
      NACK_COUNTER_TX_DMAC : out  std_logic_vector(2 downto 0);                      --! NACK counter TX
      FCT_COUNTER_TX_DMAC  : out  std_logic_vector(3 downto 0);                      --! FCT counter TX
      -- data_encapsulation (DENC) interface
      DATA_DMAC            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_encapsulation
      VALID_K_CHAR_DMAC    : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K charachter valid in the 32-bit DATA_DMAC vector
      NEW_WORD_DMAC        : out std_logic;                                          --! New word Flag to data_encapsulation
      END_PACKET_DMAC      : out std_logic;                                          --! End frame/control word to data_encapsulation
      TYPE_FRAME_DMAC      : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);   --! Type of the frame associated with DATA_DMAC
      VIRTUAL_CHANNEL_DMAC : out std_logic_vector(G_VC_NUM-1 downto 0);              --! Virtual channel of the frame associated with DATA_DMAC
      BC_TYPE_DMAC         : out std_logic_vector(G_VC_NUM-1 downto 0);              --! BROADCAST Type
      BC_CHANNEL_DMAC      : out std_logic_vector(G_VC_NUM-1 downto 0);              --! BROADCAST Channel (one channel in this implementation)
      BC_STATUS_DMAC       : out std_logic_vector(2-1 downto 0);                     --! BOADCAST status
      MULT_CHANNEL_DMAC    : out std_logic_vector(G_VC_NUM-1 downto 0);              --! Multiplier and Channel field for FCT word
      TRANS_POL_FLG_DMAC   : out std_logic;                                          --! Transmission polarity flag
      SEQ_NUM_ACK_DMAC     : out std_logic_vector(7 downto 0)                        --! SEQ_NUM ACK value
    );
  end component;

  component data_encapsulation is
    generic (
      G_VC_NUM : integer := 8                                                                     --! Number of virtual channel
    );
    port (
      CLK                               : in std_logic;                                           --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE                   : in std_logic;                                           --! Link Reset command
      -- phy_plus_lane (PPL) interface
      LANE_ACTIVE_PPL                   : in std_logic;                                           --! Lane Active flag for the DATA Link Layer
      -- data_mac (DMAC) interface
      DATA_DMAC                         : in std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel from data_mac
      VALID_K_CHAR_DMAC                 : in std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K charachter valid in the 32-bit DATA_DMAC vector
      NEW_WORD_DMAC                     : in std_logic;                                           --! New word flag from data_mac
	    END_PACKET_DMAC                   : in std_logic;                                           --! End frame/control word from data_mac
      TYPE_FRAME_DMAC                   : in std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Type of the frame associated with DATA_DMAC
      VIRTUAL_CHANNEL_DMAC              : in std_logic_vector (G_VC_NUM-1 downto 0);              --! Virtual channel of the frame associated with DATA_DMAC
      BC_TYPE_DMAC                      : in std_logic_vector (G_VC_NUM-1 downto 0);              --! BROADCAST Type
      BC_CHANNEL_DMAC                   : in std_logic_vector (G_VC_NUM-1 downto 0);              --! BROADCAST Channel (one channel in this implementation)
	    BC_STATUS_DMAC                    : in std_logic_vector (2-1 downto 0);                     --! BOADCAST status
      MULT_CHANNEL_DMAC                 : in std_logic_vector (G_VC_NUM-1 downto 0);              --! Multiplier and Channel field for FCT word
      SEQ_NUM_ACK_DMAC                  : in std_logic_vector(7 downto 0);                        --! SEQ_NUM ACK value
      TRANS_POL_FLG_DMAC                : in std_logic;                                           --! Transmission polarity flag
      -- data_seq_compute (DSCC) interface
      NEW_WORD_DENC                     : out std_logic;                                          --! New word flag to data_seq_compute
      DATA_DENC                         : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel to data_seq_compute
      VALID_K_CHARAC_DENC               : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K charachter valid in the 32-bit DATA_DENC vector
      TYPE_FRAME_DENC                   : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);   --! Type of the frame associated with DATA_DENC
      END_FRAME_DENC                    : out std_logic;                                          --! End frame/control word associated with DATA_DENC
      SEQ_NUM_ACK_DENC                  : out std_logic_vector(7 downto 0);                       --! SEQ_NUM ACK value
      TRANS_POL_FLG_DENC                : out std_logic                                           --! Transmission polarity flag
    );
  end component;

  component data_seq_compute is
    port (
	    CLK                   : in  std_logic;                                           --! Clock generated by GTY IP
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE       : in  std_logic;                                           --! Link Reset command
      -- phy_plus_lane (PPL) interface
      LANE_ACTIVE_PPL       : in  std_logic;                                           --! Lane Active flag for the DATA Link Layer
	    -- data_encapsulation (DENC) interface
	    NEW_WORD_DENC         : in  std_logic;                                           --! New word flag associated with DATA_DENC
	    DATA_DENC             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel from data_encapsulation
	    VALID_K_CHARAC_DENC   : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K charachter valid in the 32-bit DATA_DENC vector
	    TYPE_FRAME_DENC       : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Type of the frame associated with DATA_DENC
	    END_FRAME_DENC        : in  std_logic;                                           --! End frame/control word associated with DATA_DENC
	    SEQ_NUM_ACK_DENC      : in  std_logic_vector(7 downto 0);                        --! SEQ_NUM ACK value
	    TRANS_POL_FLG_DENC    : in  std_logic;                                           --! Transmission polarity flag
	    -- data_crc_compute (DCCHECK) interface
	    NEW_WORD_DSCOM        : out std_logic;                                           --! New word flag associated with DATA_DSCOM
	    DATA_DSCOM            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! Data parallel to data_encapsulation
	    VALID_K_CHARAC_DSCOM  : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! K charachter valid in the 32-bit DATA_DSCOM vector
	    TYPE_FRAME_DSCOM      : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);    --! Type of the frame associated with DATA_DSCOM
	    END_FRAME_DSCOM       : out std_logic;                                           --! End frame/control word associated with DATA_DSCOM
	    -- MIB interface
	    SEQ_NUM_DSCOM         : out std_logic_vector(7 downto 0)                         --! Current SEQ_NUM value
    );
  end component;

  component data_crc_compute is
    port (
      CLK                   : in  std_logic;                                          --! Global Clock
      -- data_link_reset (DLRE) interface
      LINK_RESET_DLRE       : in  std_logic;                                          --! Link Reset command
      -- phy_plus_lane (PPL) interface
      LANE_ACTIVE_PPL       : in  std_logic;                                          --! Lane Active flag for the DATA Link Layer
   	  -- data_seq_compute (DSCOM) interface
		  NEW_WORD_DSCOM        : in  std_logic;                                          --! New word flag associated with DATA_DSCOM
		  DATA_DSCOM            : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data parallel from data_seq_compute
		  VALID_K_CHARAC_DSCOM  : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! K charachter valid in the 32-bit DATA_DSCOM vector
		  TYPE_FRAME_DSCOM      : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);   --! Type of the frame associated with DATA_DSCOM
		  END_FRAME_DSCOM       : in  std_logic;                                          --! End frame/control word associated with DATA_DSCOM
		  -- FIFO_TX_LANE interface
		  FIFO_FULL_TX_LANE     : in  std_logic;                                          --! Fifo TX full flag from the lane layer
		  VALID_K_CHARAC_DCCOM  : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Data parallel to lane layer
		  DATA_DCCOM            : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! K charachter valid in the 32-bit DATA_DCCOM vector
		  NEW_WORD_DCCOM        : out std_logic                                           --! New word Flag associated with DATA_DCCOM
 	);
  end component;
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
  -- data_link_reset
  signal link_reset_dlre            : std_logic;
  --data_out_buf
  signal vc_ready_dobuf             : std_logic_vector(G_VC_NUM downto 0);
  signal vc_data_dobuf              : vc_data_array(G_VC_NUM downto 0);
  signal vc_valid_k_charac_dobuf    : vc_k_array(G_VC_NUM downto 0);
  signal vc_data_valid_dobuf        : std_logic_vector(G_VC_NUM downto 0);
  signal vc_end_packet_dobuf        : std_logic_vector(G_VC_NUM downto 0);
  -- data_mac
  signal req_fct_done_dmac          : std_logic_vector(G_VC_NUM-1 downto 0);
  signal req_ack_done_dmac          : std_logic;
  signal vc_rd_en_dmac              : std_logic_vector(G_VC_NUM downto 0);
  signal data_dmac                  : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dmac        : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal new_word_dmac              : std_logic;
  signal end_packet_dmac            : std_logic;
  signal type_frame_dmac            : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal virtual_channel_dmac       : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_type_dmac               : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_channel_dmac            : std_logic_vector(G_VC_NUM-1 downto 0);
  signal bc_status_dmac             : std_logic_vector(1 downto 0);
  signal mult_channel_dmac          : std_logic_vector(G_VC_NUM-1 downto 0);
  signal trans_pol_flg_dmac         : std_logic;
  signal  seq_num_ack_dmac          : std_logic_vector(7 downto 0);
  -- data_encapsulation
  signal new_word_denc              : std_logic;
  signal data_denc                  : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_denc        : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal type_frame_denc            : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal end_frame_denc             : std_logic;
  signal seq_num_ack_denc           : std_logic_vector(7 downto 0);
  signal trans_pol_flg_denc         : std_logic;
  -- data_seq_compute
  signal new_word_dscom             : std_logic;
  signal data_dscom                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dscom       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal type_frame_dscom           : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal end_frame_dscom            : std_logic;
  -- data_err_management
  signal near_end_rpf_derrm         : std_logic;
  signal req_ack_derrm              : std_logic;
  signal req_nack_derrm             : std_logic;
  signal trans_pol_flg_derrm        : std_logic;
  signal link_reset_derrm           : std_logic;
  signal  seq_num_ack_derrm         : std_logic_vector(7 downto 0);
  -- data_word_id_fsm
  signal new_word_dwi               : std_logic;
  signal end_frame_dwi              : std_logic;
  signal seq_num_dwi                : std_logic_vector(7 downto 0);
  signal crc_16b_dwi                : std_logic_vector(15 downto 0);
  signal crc_8b_dwi                 : std_logic_vector(7 downto 0);
  signal type_frame_dwi             : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal data_dwi                   : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dwi         : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal multiplier_dwi             : std_logic_vector(C_MULT_SIZE-1 downto 0);
  signal vc_dwi                     : std_logic_vector(C_CHANNEL_SIZE-1 downto 0);
  signal rxerr_dwi                  : std_logic;
  signal rxerr_all_dwi              : std_logic;
  signal frame_err_dwi              : std_logic;
  signal type_frame_dscheck         : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal rxnothing_active_dwi       : std_logic;
  -- data_crc_check
  signal seq_num_dccheck            : std_logic_vector(7 downto 0);
  signal end_frame_dccheck          : std_logic;
  signal type_frame_dccheck         : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
  signal new_word_dccheck           : std_logic;
  signal multiplier_dccheck         : std_logic_vector(C_MULT_SIZE-1 downto 0);
  signal vc_dccheck                 : std_logic_vector(C_CHANNEL_SIZE-1 downto 0);
  signal data_dccheck               : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dccheck     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal crc_err_dccheck            : std_logic;
  signal frame_err_dccheck          : std_logic;
  signal rxerr_dccheck              : std_logic;
  signal rxerr_all_dccheck          : std_logic;
  -- data_seq_check
  signal data_dscheck               : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_dscheck     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal new_word_dscheck           : std_logic;
  signal end_frame_dscheck          : std_logic;
  signal end_frame_fifo_dscheck     : std_logic;
  signal frame_err_data_dscheck     : std_logic;
  signal seq_num_err_data_dscheck   : std_logic;
  signal crc_err_data_dscheck       : std_logic;
  signal rxerr_data_dscheck         : std_logic;
  signal data_bc_dscheck            : std_logic_vector(C_DATA_LENGTH-1 downto 0);
  signal valid_k_charac_bc_dscheck  : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
  signal new_word_bc_dscheck        : std_logic;
  signal end_frame_fifo_bc_dscheck  : std_logic;
  signal frame_err_bc_dscheck       : std_logic;
  signal seq_num_err_bc_dscheck     : std_logic;
  signal crc_err_bc_dscheck         : std_logic;
  signal rxerr_bc_dscheck           : std_logic;
  signal fct_far_end_dscheck        : std_logic_vector(G_VC_NUM-1 downto 0);
  signal m_val_dscheck              : std_logic_vector(C_M_SIZE-1 downto 0);
  signal seq_num_err_dscheck        : std_logic;
  signal wr_data_dscheck            : std_logic_vector(C_DATA_K_WIDTH-1 downto 0);
  signal frame_err_dscheck          : std_logic;
  signal seq_num_ack_dscheck        : std_logic_vector(6 downto 0);
  signal crc_err_dscheck            : std_logic;
  signal rxerr_dscheck              : std_logic;
  -- data_mid_buf
  signal data_dmbuf                 : std_logic_vector(C_DATA_K_WIDTH-1 downto 0);
  signal data_rd_dmbuf              : std_logic;
  signal data_valid_dmbuf           : std_logic;
  signal status_busy_flush_dmbuf    : std_logic;
  signal frame_err_fifo_mid         : std_logic;
  -- data_desencapsulation
  signal data_ddes                  : vc_data_k_array(G_VC_NUM-1 downto 0);
  signal data_en_ddes               : std_logic_vector(G_VC_NUM-1 downto 0);
  -- data_mid_buf_bc
  signal wr_data_bc_dscheck         : std_logic_vector(C_DATA_K_WIDTH-1 downto 0);
  signal data_dmbufbc               : std_logic_vector(C_DATA_K_WIDTH-1 downto 0);
  signal data_rd_dmbufbc            : std_logic;
  signal data_valid_dmbufbc         : std_logic;
  signal status_busy_flush_dmbufbc  : std_logic;
  signal fifo_full_dmbufbc          : std_logic;
  signal frame_err_fifo_mid_bc      : std_logic;
  -- data_desencapsulation_bc
  signal data_rd_ddesbc             : std_logic;
  signal data_ddesbc                : std_logic_vector(C_DATA_K_WIDTH-1 downto 0);
  signal data_en_ddesbc             : std_logic;
  -- data_in_buf
  signal req_fct_dibuf              : std_logic_vector(G_VC_NUM-1 downto 0);
  signal link_reset_dibuf           : std_logic_vector(G_VC_NUM-1 downto 0);
begin

---------------------------------------------------------
-----                     Assignements              -----
---------------------------------------------------------
  LINK_RST_ASSERTED_DL  <= link_reset_dlre;
  SEQUENCE_ERROR_DL     <= seq_num_err_dscheck when (type_frame_dscheck /= C_ACK_FRM and type_frame_dscheck /= C_NACK_FRM) else '0';-- No sequence error for ack or nack control word
  CURRENT_TIME_SLOT_DL  <= CURRENT_TIME_SLOT_NW;
  FAR_END_LINK_RESET_DL <= FAR_END_CAPA_PPL(C_CAPA_LINK_RST);
  FRAME_ERROR_DL        <= frame_err_dwi;
  wr_data_dscheck       <= valid_k_charac_dscheck & data_dscheck;
  wr_data_bc_dscheck    <= valid_k_charac_bc_dscheck & data_bc_dscheck;
  frame_err_fifo_mid    <= seq_num_err_data_dscheck or crc_err_data_dscheck or frame_err_data_dscheck or rxerr_data_dscheck;
  frame_err_fifo_mid_bc <= seq_num_err_bc_dscheck or crc_err_bc_dscheck or frame_err_bc_dscheck or rxerr_bc_dscheck;
--------------------------------------------------------
-----                     Instantiation            -----
--------------------------------------------------------
  inst_data_in_bc_buf: data_in_bc_buf
  port map (
    RST_N                  => RST_N,
    CLK                    => CLK,
    LINK_RESET_DLRE        => link_reset_dlre,
    M_AXIS_ARSTN_NW        => AXIS_ARSTN_RX_NW(G_VC_NUM),
    M_AXIS_ACLK_NW	       => AXIS_ACLK_RX_NW(G_VC_NUM),
    M_AXIS_TVALID_DIBUF    => AXIS_TVALID_RX_DL(G_VC_NUM),
    M_AXIS_TDATA_DIBUF     => AXIS_TDATA_RX_DL(G_VC_NUM),
    M_AXIS_TLAST_DIBUF     => AXIS_TLAST_RX_DL(G_VC_NUM),
    M_AXIS_TREADY_NW       => AXIS_TREADY_RX_NW(G_VC_NUM),
    M_AXIS_TUSER_DIBUF     => AXIS_TUSER_RX_DL(G_VC_NUM),
    DATA_DDESBC            => data_ddesbc,
    DATA_EN_DDESBC         => data_en_ddesbc
  );
  inst_data_desencapsulation_bc : data_desencapsulation_bc
    port map(
      CLK                 => CLK,
      LINK_RESET_DLRE     => link_reset_dlre,
      DATA_DMBUFBC        => data_dmbufbc,
      DATA_RD_DDESBC      => data_rd_ddesbc,
      DATA_VALID_DMBUFBC  => data_valid_dmbufbc,
      DATA_DDESBC         => data_ddesbc,
      DATA_EN_DDESBC      => data_en_ddesbc
    );

  inst_mid_buf_bc: fifo_dc_drop_bad_frame
  generic map (
    G_DWIDTH            => C_DATA_K_WIDTH,
    G_AWIDTH            => C_MID_BUF_BC_SIZE
  )
  port map (
    RST_N                 => RST_N,
    WR_CLK                => CLK,
    WR_DATA               => wr_data_bc_dscheck,
    WR_DATA_EN            => new_word_bc_dscheck,
    FRAME_ERROR           => frame_err_fifo_mid_bc,
    END_FRAME             => end_frame_fifo_bc_dscheck,
    RD_CLK                => CLK,
    RD_DATA               => data_dmbufbc,
    RD_DATA_EN            => data_rd_ddesbc,
    RD_DATA_VLD           => data_valid_dmbufbc,
    CMD_FLUSH             => link_reset_dlre,
    STATUS_BUSY_FLUSH     => status_busy_flush_dmbufbc,
    STATUS_THRESHOLD_HIGH => open,
    STATUS_THRESHOLD_LOW  => open,
    STATUS_FULL           => fifo_full_dmbufbc,
    STATUS_EMPTY          => open,
    STATUS_LEVEL_WR       => open,
    STATUS_LEVEL_RD       => open
  );

  gen_data_in_buff: for i in 0 to G_VC_NUM-1 generate
    inst_data_in_buf: data_in_buf
    port map (
        RST_N                  => RST_N,
        CLK                    => CLK,
        LINK_RESET_DLRE        => link_reset_dlre,
        LINK_RESET_DIBUF       => link_reset_dibuf(i),
        M_AXIS_ARSTN_NW        => AXIS_ARSTN_RX_NW(i),
        M_AXIS_ACLK_NW	       => AXIS_ACLK_RX_NW(i),
        M_AXIS_TVALID_DIBUF    => AXIS_TVALID_RX_DL(i),
        M_AXIS_TDATA_DIBUF     => AXIS_TDATA_RX_DL(i),
        M_AXIS_TLAST_DIBUF     => AXIS_TLAST_RX_DL(i),
        M_AXIS_TREADY_NW       => AXIS_TREADY_RX_NW(i),
        M_AXIS_TUSER_DIBUF     => AXIS_TUSER_RX_DL(i),
        DATA_DDES              => data_ddes(i),
        DATA_EN_DDES           => data_en_ddes(i),
        REQ_FCT_DIBUF          => req_fct_dibuf(i),
        REQ_FCT_DONE_DMAC      => req_fct_done_dmac(i),
        INPUT_BUF_OVF_DIBUF    => INPUT_BUF_OVF_VC_DL(i)
    );
  end generate;
  inst_data_desencapsulation: data_desencapsulation
  generic map (
    G_VC_NUM => G_VC_NUM
  )
  port map (
    CLK                    => CLK,
    LINK_RESET_DLRE        => link_reset_dlre,
    DATA_DMBUF             => data_dmbuf,
    DATA_RD_DDES           => data_rd_dmbuf,
    DATA_VALID_DMBUF       => data_valid_dmbuf,
    DATA_DDES              => data_ddes,
    DATA_EN_DDES           => data_en_ddes
  );
  inst_mid_buf: fifo_dc_drop_bad_frame
  generic map (
    G_DWIDTH            => C_DATA_K_WIDTH,
    G_AWIDTH            => C_MID_BUF_SIZE
  )
  port map (
    RST_N                 => RST_N,
    WR_CLK                => CLK,
    WR_DATA               => wr_data_dscheck,
    WR_DATA_EN            => new_word_dscheck,
    FRAME_ERROR           => frame_err_fifo_mid,
    END_FRAME             => end_frame_fifo_dscheck,
    RD_CLK                => CLK,
    RD_DATA               => data_dmbuf,
    RD_DATA_EN            => data_rd_dmbuf,
    RD_DATA_VLD           => data_valid_dmbuf,
    CMD_FLUSH             => link_reset_dlre,
    STATUS_BUSY_FLUSH     => status_busy_flush_dmbuf,
    STATUS_THRESHOLD_HIGH => open,
    STATUS_THRESHOLD_LOW  => open,
    STATUS_FULL           => open,
    STATUS_EMPTY          => open,
    STATUS_LEVEL_WR       => open,
    STATUS_LEVEL_RD       => open
  );
  inst_data_seq_check: data_seq_check
  port map (
      CLK                       => CLK,
      LINK_RESET_DLRE           => link_reset_dlre,
      DATA_DCCHECK              => data_dccheck,
      VALID_K_CHARAC_DCCHECK    => valid_k_charac_dccheck,
      SEQ_NUM_DCCHECK           => seq_num_dccheck,
      END_FRAME_DCCHECK         => end_frame_dccheck,
      TYPE_FRAME_DCCHECK        => type_frame_dccheck,
      NEW_WORD_DCCHECK          => new_word_dccheck,
      CRC_ERR_DCCHECK           => crc_err_dccheck,
      FRAME_ERR_DCCHECK         => frame_err_dccheck,
      MULTIPLIER_DCCHECK        => multiplier_dccheck,
      VC_DCCHECK                => vc_dccheck,
      RXERR_DCCHECK             => rxerr_dccheck,
      RXERR_ALL_DCCHECK         => rxerr_all_dccheck,
      NEAR_END_RPF_DERRM        => near_end_rpf_derrm,
      TRANS_POL_FLG_DERRM       => trans_pol_flg_derrm,
      SEQ_NUM_ERR_DSCHECK       => seq_num_err_dscheck,
      RXERR_DSCHECK             => rxerr_dscheck,
      SEQ_NUM_ACK_DSCHECK       => seq_num_ack_dscheck,
      END_FRAME_DSCHECK         => end_frame_dscheck,
      TYPE_FRAME_DSCHECK        => type_frame_dscheck,
      DATA_DSCHECK              => data_dscheck,
      VALID_K_CHARAC_DSCHECK    => valid_k_charac_dscheck,
      NEW_WORD_DSCHECK          => new_word_dscheck,
      END_FRAME_FIFO_DSCHECK    => end_frame_fifo_dscheck,
      CRC_ERR_DSCHECK           => crc_err_dscheck,
      FRAME_ERR_DSCHECK         => frame_err_dscheck,
      FRAME_ERR_DATA_DSCHECK    => frame_err_data_dscheck,
      SEQ_NUM_ERR_DATA_DSCHECK  => seq_num_err_data_dscheck,
      CRC_ERR_DATA_DSCHECK      => crc_err_data_dscheck,
      RXERR_DATA_DSCHECK        => rxerr_data_dscheck,
      DATA_BC_DSCHECK           => data_bc_dscheck,
      VALID_K_CHARAC_BC_DSCHECK => valid_k_charac_bc_dscheck,
      NEW_WORD_BC_DSCHECK       => new_word_bc_dscheck,
      END_FRAME_FIFO_BC_DSCHECK => end_frame_fifo_bc_dscheck,
      FRAME_ERR_BC_DSCHECK      => frame_err_bc_dscheck,
      SEQ_NUM_ERR_BC_DSCHECK    => seq_num_err_bc_dscheck,
      CRC_ERR_BC_DSCHECK        => crc_err_bc_dscheck,
      RXERR_BC_DSCHECK          => rxerr_bc_dscheck,
      FCT_FAR_END_DSCHECK       => fct_far_end_dscheck,
      M_VAL_DSCHECK             => m_val_dscheck,
      SEQ_NUM_DSCHECK           => SEQ_NUMBER_RX_DL,
      NACK_SEQ_NUM_DSCHECK      => NACK_SEQ_NUM_DL,
      ACK_SEQ_NUM_DSCHECK       => ACK_SEQ_NUM_DL,
      ACK_COUNTER_RX_DSCHECK    => ACK_COUNTER_RX_DL,
      NACK_COUNTER_RX_DSCHECK   => NACK_COUNTER_RX_DL,
      FCT_COUNTER_RX_DSCHECK    => FCT_COUNTER_RX_DL,
      FULL_COUNTER_RX_DSCHECK   => FULL_COUNTER_RX_DL,
      ACK_PULSE_RX_DSCHECK      => ACK_PULSE_RX_DL,
      NACK_PULSE_RX_DSCHECK     => NACK_PULSE_RX_DL,
      FCT_PULSE_RX_DSCHECK      => FCT_PULSE_RX_DL,
      FULL_PULSE_RX_DSCHECK     => FULL_PULSE_RX_DL
  );

  inst_data_crc_check: data_crc_check
  port map (
      CLK                    => CLK,
      LINK_RESET_DLRE        => link_reset_dlre,
      DATA_DWI               => data_dwi,
      VALID_K_CHARAC_DWI     => valid_k_charac_dwi,
      NEW_WORD_DWI           => new_word_dwi,
      END_FRAME_DWI          => end_frame_dwi,
      SEQ_NUM_DWI            => seq_num_dwi,
      CRC_16B_DWI            => crc_16b_dwi,
      CRC_8B_DWI             => crc_8b_dwi,
      MULTIPLIER_DWI         => multiplier_dwi,
      VC_DWI                 => vc_dwi,
      TYPE_FRAME_DWI         => type_frame_dwi,
      FRAME_ERR_DWI          => frame_err_dwi,
      RXERR_DWI              => rxerr_dwi,
      RXERR_ALL_DWI           => rxerr_all_dwi,
      RXNOTHING_ACTIVE_DWI   => rxnothing_active_dwi,
      NEW_WORD_DCCHECK       => new_word_dccheck,
      DATA_DCCHECK           => data_dccheck,
      VALID_K_CHARAC_DCCHECK => valid_k_charac_dccheck,
      END_FRAME_DCCHECK      => end_frame_dccheck,
      TYPE_FRAME_DCCHECK     => type_frame_dccheck,
      SEQ_NUM_DCCHECK        => seq_num_dccheck,
      CRC_ERR_DCCHECK        => crc_err_dccheck,
      FRAME_ERR_DCCHECK      => frame_err_dccheck,
      MULTIPLIER_DCCHECK     => multiplier_dccheck,
      VC_DCCHECK             => vc_dccheck,
      RXERR_DCCHECK          => rxerr_dccheck,
      RXERR_ALL_DCCHECK      => rxerr_all_dccheck,
      CRC_LONG_ERR_DCCHECK   => CRC_LONG_ERROR_DL,
      CRC_SHORT_ERR_DCCHECK  => CRC_SHORT_ERROR_DL
  );
  inst_data_word_id_fsm: data_word_id_fsm
  port map (
      CLK                     => CLK,
      LINK_RESET_DLRE         => link_reset_dlre,
      FIFO_RX_DATA_VALID_PPL  => FIFO_RX_DATA_VALID_PPL,
      FIFO_RX_RD_EN_DL        => FIFO_RX_RD_EN_DL,
      DATA_RX_PPL             => DATA_RX_PPL,
      VALID_K_CHARAC_PPL      => VALID_K_CHARAC_RX_PPL,
      TYPE_FRAME_DWI          => type_frame_dwi,
      NEW_WORD_DWI            => new_word_dwi,
      END_FRAME_DWI           => end_frame_dwi,
      DATA_DWI                => data_dwi,
      VALID_K_CHARAC_DWI      => valid_k_charac_dwi,
      SEQ_NUM_DWI             => seq_num_dwi,
      CRC_16B_DWI             => crc_16b_dwi,
      CRC_8B_DWI              => crc_8b_dwi,
      MULTIPLIER_DWI          => multiplier_dwi,
      VC_DWI                  => vc_dwi,
      RXNOTHING_ACTIVE_DWI    => rxnothing_active_dwi,
      CRC_ERR_DCCHECK         => crc_err_dccheck,
      SEQ_ERR_DSCHECK         => seq_num_err_dscheck,
      FRAME_ERR_DWI           => frame_err_dwi,
      RXERR_DWI               => rxerr_dwi,
      RXERR_ALL_DWI           => rxerr_all_dwi,
      DATA_COUNTER_RX_DWI     => DATA_COUNTER_RX_DL,
      RETRY_COUNTER_RX_DWI    => RETRY_COUNTER_RX_DL,
      DATA_PULSE_RX_DWI       => DATA_PULSE_RX_DL,
      RETRY_PULSE_RX_DWI      => RETRY_PULSE_RX_DL
  );
  inst_data_err_management: data_err_management
  port map (
      CLK                      => CLK,
      LINK_RESET_DLRE          => link_reset_dlre,
      LINK_RESET_DERRM         => link_reset_derrm,
      RXERR_DSCHECK            => rxerr_dscheck,
      CRC_ERR_DSCHECK          => crc_err_dscheck,
      TYPE_FRAME_DSCHECK       => type_frame_dscheck,
      END_FRAME_DSCHECK        => end_frame_dscheck,
      SEQ_ERR_DSCHECK          => seq_num_err_dscheck,
      SEQ_NUM_ACK_DSCHECK      => seq_num_ack_dscheck,
      FAR_END_RPF_DSCHECK      => '0',
      NEAR_END_RPF_DERRM       => near_end_rpf_derrm,
      FRAME_ERR_DSCHECK        => frame_err_dscheck,
      REQ_ACK_DERRM            => req_ack_derrm,
      REQ_NACK_DERRM           => req_nack_derrm,
      TRANS_POL_FLG_DERRM      => trans_pol_flg_derrm,
      SEQ_NUM_ACK_DERRM        => seq_num_ack_derrm,
      REQ_ACK_DONE_DMAC        => req_ack_done_dmac,
      NACK_RST_EN_MIB          => NACK_RST_EN_MIB,
      NACK_RST_MODE_MIB        => NACK_RST_MODE_MIB
  );
  inst_data_link_reset: data_link_reset
  generic map (
    G_VC_NUM => G_VC_NUM
  )
  port map (
      RST_N                   => RST_N,
      CLK                     => CLK,
      LINK_RESET_DLRE         => link_reset_dlre,
      LINK_RESET_DIBUF        => link_reset_dibuf,
      LINK_RESET_DERRM        => link_reset_derrm,
      RESET_PARAM_DLRE        => RESET_PARAM_DL,
      LANE_RESET_DLRE         => LANE_RESET_DL,
      NEAR_END_CAPA_DLRE      => CAPABILITY_TX_DL,
      LANE_ACTIVE_PPL         => LANE_ACTIVE_PPL,
      FAR_END_CAPA_PPL        => FAR_END_CAPA_PPL,
      INTERFACE_RESET_MIB     => INTERFACE_RESET_MIB,
      LINK_RESET_MIB          => LINK_RESET_MIB
  );
  inst_data_out_bc_buf: data_out_bc_buf
    port map (
      RST_N                 => RST_N,
      CLK                   => CLK,
      LINK_RESET_DLRE       => link_reset_dlre,
      S_AXIS_ARSTN_NW       => AXIS_ARSTN_TX_NW(G_VC_NUM),
      S_AXIS_ACLK_NW	    => AXIS_ACLK_TX_NW(G_VC_NUM),
      S_AXIS_TREADY_DL      => AXIS_TREADY_TX_DL(G_VC_NUM),
      S_AXIS_TDATA_NW       => AXIS_TDATA_TX_NW(G_VC_NUM),
      S_AXIS_TUSER_NW       => AXIS_TUSER_TX_NW(G_VC_NUM),
      S_AXIS_TLAST_NW       => AXIS_TLAST_TX_NW(G_VC_NUM),
      S_AXIS_TVALID_NW      => AXIS_TVALID_TX_NW(G_VC_NUM),
      VC_READY_DOBUF        => vc_ready_dobuf(G_VC_NUM),
      DATA_DOBUF            => vc_data_dobuf(G_VC_NUM),
      VALID_K_CHARAC_DOBUF  => vc_valid_k_charac_dobuf(G_VC_NUM),
      DATA_VALID_DOBUF      => vc_data_valid_dobuf(G_VC_NUM),
      END_PACKET_DOBUF      => vc_end_packet_dobuf(G_VC_NUM),
      VC_RD_EN_DMAC         => vc_rd_en_dmac(G_VC_NUM)
    );
 
  gen_data_out_buff: for i in 0 to G_VC_NUM-1 generate
    inst_data_out_buff: data_out_buff
      port map (
        RST_N                 => RST_N,
        CLK                   => CLK,
        LINK_RESET_DLRE       => link_reset_dlre,
        S_AXIS_ARSTN_NW       => AXIS_ARSTN_TX_NW(i),
        S_AXIS_ACLK_NW	      => AXIS_ACLK_TX_NW(i),
        S_AXIS_TREADY_DL      => AXIS_TREADY_TX_DL(i),
        S_AXIS_TDATA_NW       => AXIS_TDATA_TX_NW(i),
        S_AXIS_TUSER_NW       => AXIS_TUSER_TX_NW(i),
        S_AXIS_TLAST_NW       => AXIS_TLAST_TX_NW(i),
        S_AXIS_TVALID_NW      => AXIS_TVALID_TX_NW(i),
        VC_READY_DOBUF        => vc_ready_dobuf(i),
        DATA_DOBUF            => vc_data_dobuf(i),
        VALID_K_CHARAC_DOBUF  => vc_valid_k_charac_dobuf(i),
        DATA_VALID_DOBUF      => vc_data_valid_dobuf(i),
        END_PACKET_DOBUF      => vc_end_packet_dobuf(i),
        VC_RD_EN_DMAC         => vc_rd_en_dmac(i),
        M_VAL_DSCHECK         => m_val_dscheck,
        FCT_FAR_END_DSCHECK   => fct_far_end_dscheck(i),
        LANE_ACTIVE_ST_PPL    => LANE_ACTIVE_PPL,
        FCT_CC_OVF_DOBUF      => FCT_CREDIT_OVERFLOW_DL(i),
        CREDIT_VC_DOBUF       => CREDIT_VC_DL(i),
        VC_CONT_MODE_MIB      => CONTINUOUS_VC_MIB(i)
      );
  end generate;
  inst_data_mac: data_mac
    generic map (
      G_VC_NUM => G_VC_NUM
    )
    port map (
      CLK                  => CLK,
      LINK_RESET_DLRE      => link_reset_dlre,
      LANE_ACTIVE_PPL      => LANE_ACTIVE_PPL,
      REQ_ACK_DERRM        => req_ack_derrm,
      REQ_NACK_DERRM       => req_nack_derrm,
      TRANS_POL_FLG_DERRM  => trans_pol_flg_derrm,
      REQ_ACK_DONE_DMAC    => req_ack_done_dmac,
      SEQ_NUM_ACK_DERRM    => seq_num_ack_derrm,
      REQ_FCT_DONE_DMAC    => req_fct_done_dmac,
      REQ_FCT_DIBUF        => req_fct_dibuf,
      VC_READY_DOBUF       => vc_ready_dobuf,
      VC_DATA_DOBUF        => vc_data_dobuf,
      VC_VALID_K_CHAR_DOBUF=> vc_valid_k_charac_dobuf,
      VC_DATA_VALID_DOBUF  => vc_data_valid_dobuf,
      VC_END_PACKET_DOBUF  => vc_end_packet_dobuf,
      VC_RD_EN_DMAC        => vc_rd_en_dmac,
      VC_PAUSE_MIB         => PAUSE_VC_MIB,
      VC_END_EMISSION_DMAC => FRAME_FINISHED_DL,
      VC_RUN_EMISSION_DMAC => FRAME_TX_DL,
      DATA_COUNTER_TX_DMAC => DATA_COUNTER_TX_DL,
      ACK_COUNTER_TX_DMAC  => ACK_COUNTER_TX_DL,
      NACK_COUNTER_TX_DMAC => NACK_COUNTER_TX_DL,
      FCT_COUNTER_TX_DMAC  => FCT_COUNTER_TX_DL,
      DATA_DMAC            => data_dmac,
      VALID_K_CHAR_DMAC    => valid_k_charac_dmac,
      NEW_WORD_DMAC        => new_word_dmac,
      END_PACKET_DMAC      => end_packet_dmac,
      TYPE_FRAME_DMAC      => type_frame_dmac,
      VIRTUAL_CHANNEL_DMAC => virtual_channel_dmac,
      BC_TYPE_DMAC         => bc_type_dmac,
      BC_CHANNEL_DMAC      => bc_channel_dmac,
      BC_STATUS_DMAC       => bc_status_dmac,
      MULT_CHANNEL_DMAC    => mult_channel_dmac,
      TRANS_POL_FLG_DMAC   => trans_pol_flg_dmac,
      SEQ_NUM_ACK_DMAC     => seq_num_ack_dmac
    );

  inst_data_encapsulation: data_encapsulation
    generic map (
      G_VC_NUM => G_VC_NUM
    )
    port map (
      CLK                   => CLK,
      LINK_RESET_DLRE       => link_reset_dlre,
      LANE_ACTIVE_PPL       => LANE_ACTIVE_PPL,
      DATA_DMAC             => data_dmac,
      VALID_K_CHAR_DMAC     => valid_k_charac_dmac,
      NEW_WORD_DMAC         => new_word_dmac,
      END_PACKET_DMAC       => end_packet_dmac,
      TYPE_FRAME_DMAC       => type_frame_dmac,
      VIRTUAL_CHANNEL_DMAC  => virtual_channel_dmac,
      BC_TYPE_DMAC          => bc_type_dmac,
      BC_CHANNEL_DMAC       => bc_channel_dmac,
      BC_STATUS_DMAC        => bc_status_dmac,
      MULT_CHANNEL_DMAC     => mult_channel_dmac,
      SEQ_NUM_ACK_DMAC      => seq_num_ack_dmac,
      TRANS_POL_FLG_DMAC    => trans_pol_flg_dmac,
      NEW_WORD_DENC         => new_word_denc,
      DATA_DENC             => data_denc,
      VALID_K_CHARAC_DENC   => valid_k_charac_denc,
      TYPE_FRAME_DENC       => type_frame_denc,
      END_FRAME_DENC        => end_frame_denc,
      SEQ_NUM_ACK_DENC      => seq_num_ack_denc,
      TRANS_POL_FLG_DENC    => trans_pol_flg_denc
    );

  inst_data_seq_compute: data_seq_compute
    port map (
      CLK                   => CLK,
      LINK_RESET_DLRE       => link_reset_dlre,
      LANE_ACTIVE_PPL       => LANE_ACTIVE_PPL,
      NEW_WORD_DENC         => new_word_denc,
      DATA_DENC             => data_denc,
      VALID_K_CHARAC_DENC   => valid_k_charac_denc,
      TYPE_FRAME_DENC       => type_frame_denc,
      END_FRAME_DENC        => end_frame_denc,
      SEQ_NUM_ACK_DENC      => seq_num_ack_denc,
      TRANS_POL_FLG_DENC    => trans_pol_flg_denc,
      NEW_WORD_DSCOM        => new_word_dscom,
      DATA_DSCOM            => data_dscom,
      VALID_K_CHARAC_DSCOM  => valid_k_charac_dscom,
      TYPE_FRAME_DSCOM      => type_frame_dscom,
      END_FRAME_DSCOM       => end_frame_dscom,
      SEQ_NUM_DSCOM         => SEQ_NUMBER_TX_DL
    );

  inst_data_crc_compute: data_crc_compute
    port map (
      CLK                   => CLK,
      LINK_RESET_DLRE       => link_reset_dlre,
      LANE_ACTIVE_PPL       => LANE_ACTIVE_PPL,
      NEW_WORD_DSCOM        => new_word_dscom,
      DATA_DSCOM            => data_dscom,
      VALID_K_CHARAC_DSCOM  => valid_k_charac_dscom,
      TYPE_FRAME_DSCOM      => type_frame_dscom,
      END_FRAME_DSCOM       => end_frame_dscom,
      FIFO_FULL_TX_LANE     => FIFO_TX_FULL_PPL,
      VALID_K_CHARAC_DCCOM  => VALID_K_CHARAC_TX_DL,
      DATA_DCCOM            => DATA_TX_DL,
      NEW_WORD_DCCOM        => NEW_DATA_TX_DL
    );
end Behavioral;
