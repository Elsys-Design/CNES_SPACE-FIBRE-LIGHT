// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_RAM32X16DR8_DEFINES_VH
`else
`define B_RAM32X16DR8_DEFINES_VH

// Look-up table parameters
//

`define RAM32X16DR8_ADDR_N  9
`define RAM32X16DR8_ADDR_SZ 32
`define RAM32X16DR8_DATA_SZ 64

// Attribute addresses
//

`define RAM32X16DR8__INIT_A    32'h00000000
`define RAM32X16DR8__INIT_A_SZ 64

`define RAM32X16DR8__INIT_B    32'h00000001
`define RAM32X16DR8__INIT_B_SZ 64

`define RAM32X16DR8__INIT_C    32'h00000002
`define RAM32X16DR8__INIT_C_SZ 64

`define RAM32X16DR8__INIT_D    32'h00000003
`define RAM32X16DR8__INIT_D_SZ 64

`define RAM32X16DR8__INIT_E    32'h00000004
`define RAM32X16DR8__INIT_E_SZ 64

`define RAM32X16DR8__INIT_F    32'h00000005
`define RAM32X16DR8__INIT_F_SZ 64

`define RAM32X16DR8__INIT_G    32'h00000006
`define RAM32X16DR8__INIT_G_SZ 64

`define RAM32X16DR8__INIT_H    32'h00000007
`define RAM32X16DR8__INIT_H_SZ 64

`define RAM32X16DR8__IS_WCLK_INVERTED    32'h00000008
`define RAM32X16DR8__IS_WCLK_INVERTED_SZ 1

`endif  // B_RAM32X16DR8_DEFINES_VH