`include "B_IDELAYE3_defines.vh"

reg [`IDELAYE3_DATA_SZ-1:0] ATTR [0:`IDELAYE3_ADDR_N-1];
reg [`IDELAYE3__CASCADE_SZ:1] CASCADE_REG = CASCADE;
reg [`IDELAYE3__DELAY_FORMAT_SZ:1] DELAY_FORMAT_REG = DELAY_FORMAT;
reg [`IDELAYE3__DELAY_SRC_SZ:1] DELAY_SRC_REG = DELAY_SRC;
reg [`IDELAYE3__DELAY_TYPE_SZ:1] DELAY_TYPE_REG = DELAY_TYPE;
reg [`IDELAYE3__DELAY_VALUE_SZ-1:0] DELAY_VALUE_REG = DELAY_VALUE;
reg IS_CLK_INVERTED_REG = IS_CLK_INVERTED;
reg IS_RST_INVERTED_REG = IS_RST_INVERTED;
reg [`IDELAYE3__LOOPBACK_SZ:1] LOOPBACK_REG = LOOPBACK;
real REFCLK_FREQUENCY_REG = REFCLK_FREQUENCY;
reg [`IDELAYE3__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
real SIM_VERSION_REG = SIM_VERSION;
reg [`IDELAYE3__UPDATE_MODE_SZ:1] UPDATE_MODE_REG = UPDATE_MODE;

initial begin
  ATTR[`IDELAYE3__CASCADE] = CASCADE;
  ATTR[`IDELAYE3__DELAY_FORMAT] = DELAY_FORMAT;
  ATTR[`IDELAYE3__DELAY_SRC] = DELAY_SRC;
  ATTR[`IDELAYE3__DELAY_TYPE] = DELAY_TYPE;
  ATTR[`IDELAYE3__DELAY_VALUE] = DELAY_VALUE;
  ATTR[`IDELAYE3__IS_CLK_INVERTED] = IS_CLK_INVERTED;
  ATTR[`IDELAYE3__IS_RST_INVERTED] = IS_RST_INVERTED;
  ATTR[`IDELAYE3__LOOPBACK] = LOOPBACK;
  ATTR[`IDELAYE3__REFCLK_FREQUENCY] = $realtobits(REFCLK_FREQUENCY);
  ATTR[`IDELAYE3__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`IDELAYE3__SIM_VERSION] = $realtobits(SIM_VERSION);
  ATTR[`IDELAYE3__UPDATE_MODE] = UPDATE_MODE;
end

always @(trig_attr) begin
  CASCADE_REG = ATTR[`IDELAYE3__CASCADE];
  DELAY_FORMAT_REG = ATTR[`IDELAYE3__DELAY_FORMAT];
  DELAY_SRC_REG = ATTR[`IDELAYE3__DELAY_SRC];
  DELAY_TYPE_REG = ATTR[`IDELAYE3__DELAY_TYPE];
  DELAY_VALUE_REG = ATTR[`IDELAYE3__DELAY_VALUE];
  IS_CLK_INVERTED_REG = ATTR[`IDELAYE3__IS_CLK_INVERTED];
  IS_RST_INVERTED_REG = ATTR[`IDELAYE3__IS_RST_INVERTED];
  LOOPBACK_REG = ATTR[`IDELAYE3__LOOPBACK];
  REFCLK_FREQUENCY_REG = $bitstoreal(ATTR[`IDELAYE3__REFCLK_FREQUENCY]);
  SIM_DEVICE_REG = ATTR[`IDELAYE3__SIM_DEVICE];
  SIM_VERSION_REG = $bitstoreal(ATTR[`IDELAYE3__SIM_VERSION]);
  UPDATE_MODE_REG = ATTR[`IDELAYE3__UPDATE_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IDELAYE3_ADDR_SZ-1:0] addr;
  input  [`IDELAYE3_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IDELAYE3_DATA_SZ-1:0] read_attr;
  input  [`IDELAYE3_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
