`include "B_DSP_FP_OUTPUT_TEST_defines.vh"

reg [`DSP_FP_OUTPUT_TEST_DATA_SZ-1:0] ATTR [0:`DSP_FP_OUTPUT_TEST_ADDR_N-1];
reg [56:1] EN_SCAN_REG = EN_SCAN;
reg [31:0] FPA_PREG_REG = FPA_PREG;
reg [31:0] FPM_PREG_REG = FPM_PREG;
reg IS_RSTFPA_INVERTED_REG = IS_RSTFPA_INVERTED;
reg IS_RSTFPM_INVERTED_REG = IS_RSTFPM_INVERTED;
reg [40:1] LEGACY_REG = LEGACY;
reg [24:1] PCOUTSEL_REG = PCOUTSEL;
reg [40:1] RESET_MODE_REG = RESET_MODE;
reg [64:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_FP_OUTPUT_TEST__EN_SCAN] = EN_SCAN;
  ATTR[`DSP_FP_OUTPUT_TEST__FPA_PREG] = FPA_PREG;
  ATTR[`DSP_FP_OUTPUT_TEST__FPM_PREG] = FPM_PREG;
  ATTR[`DSP_FP_OUTPUT_TEST__IS_RSTFPA_INVERTED] = IS_RSTFPA_INVERTED;
  ATTR[`DSP_FP_OUTPUT_TEST__IS_RSTFPM_INVERTED] = IS_RSTFPM_INVERTED;
  ATTR[`DSP_FP_OUTPUT_TEST__LEGACY] = LEGACY;
  ATTR[`DSP_FP_OUTPUT_TEST__PCOUTSEL] = PCOUTSEL;
  ATTR[`DSP_FP_OUTPUT_TEST__RESET_MODE] = RESET_MODE;
  ATTR[`DSP_FP_OUTPUT_TEST__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  EN_SCAN_REG = ATTR[`DSP_FP_OUTPUT_TEST__EN_SCAN];
  FPA_PREG_REG = ATTR[`DSP_FP_OUTPUT_TEST__FPA_PREG];
  FPM_PREG_REG = ATTR[`DSP_FP_OUTPUT_TEST__FPM_PREG];
  IS_RSTFPA_INVERTED_REG = ATTR[`DSP_FP_OUTPUT_TEST__IS_RSTFPA_INVERTED];
  IS_RSTFPM_INVERTED_REG = ATTR[`DSP_FP_OUTPUT_TEST__IS_RSTFPM_INVERTED];
  LEGACY_REG = ATTR[`DSP_FP_OUTPUT_TEST__LEGACY];
  PCOUTSEL_REG = ATTR[`DSP_FP_OUTPUT_TEST__PCOUTSEL];
  RESET_MODE_REG = ATTR[`DSP_FP_OUTPUT_TEST__RESET_MODE];
  USE_MULT_REG = ATTR[`DSP_FP_OUTPUT_TEST__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_FP_OUTPUT_TEST_ADDR_SZ-1:0] addr;
  input  [`DSP_FP_OUTPUT_TEST_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_FP_OUTPUT_TEST_DATA_SZ-1:0] read_attr;
  input  [`DSP_FP_OUTPUT_TEST_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
