// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_CPM5N_DEFINES_VH
`else
`define B_CPM5N_DEFINES_VH

// Look-up table parameters
//

`define CPM5N_ADDR_N  19
`define CPM5N_ADDR_SZ 32
`define CPM5N_DATA_SZ 184

// Attribute addresses
//

`define CPM5N__CDX_MODE    32'h00000000
`define CPM5N__CDX_MODE_SZ 32

`define CPM5N__CPM5N_MPIOBOT_MODE    32'h00000001
`define CPM5N__CPM5N_MPIOBOT_MODE_SZ 160

`define CPM5N__CPM5N_MPIOTOP_MODE    32'h00000002
`define CPM5N__CPM5N_MPIOTOP_MODE_SZ 160

`define CPM5N__DPU_MODE    32'h00000003
`define CPM5N__DPU_MODE_SZ 80

`define CPM5N__LINK_SPEED_0    32'h00000004
`define CPM5N__LINK_SPEED_0_SZ 48

`define CPM5N__LINK_SPEED_1    32'h00000005
`define CPM5N__LINK_SPEED_1_SZ 32

`define CPM5N__LINK_SPEED_2    32'h00000006
`define CPM5N__LINK_SPEED_2_SZ 48

`define CPM5N__LINK_SPEED_3    32'h00000007
`define CPM5N__LINK_SPEED_3_SZ 32

`define CPM5N__LINK_WIDTH_0    32'h00000008
`define CPM5N__LINK_WIDTH_0_SZ 5

`define CPM5N__LINK_WIDTH_1    32'h00000009
`define CPM5N__LINK_WIDTH_1_SZ 3

`define CPM5N__LINK_WIDTH_2    32'h0000000a
`define CPM5N__LINK_WIDTH_2_SZ 4

`define CPM5N__LINK_WIDTH_3    32'h0000000b
`define CPM5N__LINK_WIDTH_3_SZ 3

`define CPM5N__PACKET_SIZE    32'h0000000c
`define CPM5N__PACKET_SIZE_SZ 11

`define CPM5N__PCIE_MODE_A0    32'h0000000d
`define CPM5N__PCIE_MODE_A0_SZ 184

`define CPM5N__PCIE_MODE_A1    32'h0000000e
`define CPM5N__PCIE_MODE_A1_SZ 184

`define CPM5N__PCIE_MODE_A2    32'h0000000f
`define CPM5N__PCIE_MODE_A2_SZ 184

`define CPM5N__PCIE_MODE_A3    32'h00000010
`define CPM5N__PCIE_MODE_A3_SZ 184

`define CPM5N__SIM_CPM_CDO_FILE_NAME    32'h00000011
`define CPM5N__SIM_CPM_CDO_FILE_NAME_SZ 88

`define CPM5N__SIM_CPM_CDO_MODE    32'h00000012
`define CPM5N__SIM_CPM_CDO_MODE_SZ 2

`endif  // B_CPM5N_DEFINES_VH