// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IBUFDS_INTERMDISABLE_DEFINES_VH
`else
`define B_IBUFDS_INTERMDISABLE_DEFINES_VH

// Look-up table parameters
//

`define IBUFDS_INTERMDISABLE_ADDR_N  6
`define IBUFDS_INTERMDISABLE_ADDR_SZ 32
`define IBUFDS_INTERMDISABLE_DATA_SZ 88

// Attribute addresses
//

`define IBUFDS_INTERMDISABLE__DIFF_TERM    32'h00000000
`define IBUFDS_INTERMDISABLE__DIFF_TERM_SZ 40

`define IBUFDS_INTERMDISABLE__DQS_BIAS    32'h00000001
`define IBUFDS_INTERMDISABLE__DQS_BIAS_SZ 40

`define IBUFDS_INTERMDISABLE__IBUF_LOW_PWR    32'h00000002
`define IBUFDS_INTERMDISABLE__IBUF_LOW_PWR_SZ 40

`define IBUFDS_INTERMDISABLE__IOSTANDARD    32'h00000003
`define IBUFDS_INTERMDISABLE__IOSTANDARD_SZ 56

`define IBUFDS_INTERMDISABLE__SIM_DEVICE    32'h00000004
`define IBUFDS_INTERMDISABLE__SIM_DEVICE_SZ 88

`define IBUFDS_INTERMDISABLE__USE_IBUFDISABLE    32'h00000005
`define IBUFDS_INTERMDISABLE__USE_IBUFDISABLE_SZ 40

`endif  // B_IBUFDS_INTERMDISABLE_DEFINES_VH