-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
--------------------------------------------------------------------------
-- COMPANY       : CNES
--------------------------------------------------------------------------
-- TITLE         : data_link_configurator.vhd
-- PROJECT       : SPACE FIBRE LIGHT
--------------------------------------------------------------------------
-- AUTHOR        : Thomas Favre Felix
-- CREATED       : 12/03/2024
--------------------------------------------------------------------------
-- DESCRIPTION   : Model able to communicate with IP PHY/LANE/DATA LINK
--                 MIB blocks
--------------------------------------------------------------------------
-- History       : V1.0: Creation of the file
--------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_model.all;
------------------------------------------------------------------------------------------------------------------
--                                                      ENTITY                                                  --
------------------------------------------------------------------------------------------------------------------
entity DATA_LINK_CONFIGURATOR is
    generic(
       G_ADDR_WIDTH : positive := C_AXI_ADDR_WIDTH;                              -- Generic for AXI address width
       G_DATA_WIDTH : positive := C_AXI_DATA_WIDTH;                              -- Generic for AXI data width
       G_CHANNEL_NUMBER : positive := C_CHANNEL_NUMBER                           -- Generic for number of channel
    );
    port(
   -- Clock and reset
   ------------------
   CLK                   : in std_logic;                                         -- Clock signal
   RST_N                 : in std_logic;                                         -- Reset active low signal
   CLK_TX                : in  std_logic;                                        -- Clock generated by manufacturer IP
   RST_TXCLK_N           : in  std_logic;                                        -- Reset clock generated by manufacturer IP
   CLK_DL                : in  std_logic;                                        -- Clock of the Data Link layer
   RST_N_DL              : in std_logic;                                         -- Reset active low signal from Data Link layer
   -- AXI4 Lite slave interface
   ---------------------------------------
       -- Write Address channel (AW)
   S_AXI_AWADDR          : in std_logic_vector(G_ADDR_WIDTH-1 downto 0);         -- Write address from master to slave
   S_AXI_AWVALID         : in std_logic;                                         -- Master asserts when write address is valid
   S_AXI_AWREADY         : out std_logic;                                        -- Slave ready to accept write address
       -- Write Data channel (W)
   S_AXI_WDATA           : in std_logic_vector(G_DATA_WIDTH-1 downto 0);         -- Write data from master
   S_AXI_WSTRB           : in std_logic_vector(3 downto 0);                      -- Write strobe, indicates active byte lanes
   S_AXI_WVALID          : in std_logic;                                         -- Master asserts when write data is valid
   S_AXI_WREADY          : out std_logic;                                        -- Slave ready to accept write data
       -- Write Response channel (B)
   S_AXI_BREADY          : in std_logic;                                         -- Master ready to receive write response
   S_AXI_BRESP           : out std_logic_vector(1 downto 0);                     -- Write response from slave (OKAY or ERROR)
   S_AXI_BVALID          : out std_logic;                                        -- Slave asserts when write response is valid
       --Read Address channel (AR)
   S_AXI_ARADDR          : in std_logic_vector(G_ADDR_WIDTH-1 downto 0);         -- Read address from master to slave
   S_AXI_ARVALID         : in std_logic;                                         -- Master asserts when read address is valid
   S_AXI_ARREADY         : out std_logic;                                        -- Slave ready to accept read address
       -- Read channel (R)
   S_AXI_RREADY          : in std_logic;                                         -- Master ready to receive read data
   S_AXI_RDATA           : out std_logic_vector(G_DATA_WIDTH-1 downto 0);        -- Read data from slave to master
   S_AXI_RRESP           : out std_logic_vector(1 downto 0);                     -- Read response (OKAY or ERROR)
   S_AXI_RVALID          : out std_logic;                                        -- Slave asserts when read data is valid

   -- LANE + PHY interface
   ---------------------------------------
   -- to the DATA LINK
   INTERFACE_RST         : out std_logic;                                        -- Enable interface reset
   LINK_RST              : out std_logic;                                        -- Reset link
   NACK_RST_EN           : out std_logic;                                        -- Enable automatic reset on NACK reception
   NACK_RST_MODE         : out std_logic;                                        -- Select automatic reset mode on NACK reception
   PAUSE_VC              : out std_logic_vector(G_CHANNEL_NUMBER downto 0);      -- Pause each corresponding channel at the end of the current frame being sent
   CONTINUOUS_VC         : out std_logic_vector(G_CHANNEL_NUMBER-1 downto 0);    -- Enable continuous mode of each corresponding virtual channel

   -- to the LANE
   LANE_START            : out std_logic;                                        -- SpaceFibre lane start initialization signal
   AUTOSTART             : out std_logic;                                        -- Enables communication lane to initialize automatically when a link is established
   LANE_RESET            : out std_logic;                                        -- Reset Lane layer signal
   PARALLEL_LOOPBACK_EN  : out std_logic;                                        -- Parallel loopback enables signal
   STANDBY_REASON        : out std_logic_vector(C_STDBYREASON_WIDTH-1 downto 0); -- Standby reason field

   -- to the PHY
   NEAR_END_SERIAL_LB_EN : out std_logic;                                        -- Near-End Serial Loopback
   FAR_END_SERIAL_LB_EN  : out std_logic;                                        -- Far -End Serial Loopback

   -- from the DATA LINK
   VC_CREDIT             : in std_logic_vector(G_CHANNEL_NUMBER-1 downto 0);     -- Up if each corresponding virtual channel has credit in the far-end input buffer
   FCT_CREDIT_OVERFLOW   : in std_logic_vector(G_CHANNEL_NUMBER-1 downto 0);     -- Up if each corresponding virtual channel credit counter overflowed
   CRC_LONG_ERROR        : in std_logic;                                         -- RX error in CRC-16bit
   CRC_SHORT_ERROR       : in std_logic;                                         -- RX error in CRC-8bit
   FRAME_ERROR           : in std_logic;                                         -- RX frame error
   SEQ_ERROR             : in std_logic;                                         -- RX SEQUENCE_NUMBER error
   FAR_END_LINK_RST      : in std_logic;                                         -- Far-end Link reset status
   SEQ_NUMBER_TX         : in std_logic_vector(7 downto 0);                      -- SEQ_NUMBER in transmission
   SEQ_NUMBER_RX         : in std_logic_vector(7 downto 0);                      -- SEQ_NUMBER in reception
   INPUT_BUFFER_OVFL     : in std_logic_vector(7 downto 0);                      -- Up if the corresponding input buffer has overflowed
   FRAME_TX              : in std_logic_vector(8 downto 0);
   FRAME_FINISHED        : in std_logic_vector(8 downto 0);
   DATA_CNT_TX           : in std_logic_vector(6 downto 0);
   DATA_CNT_RX           : in std_logic_vector(6 downto 0);
   ACK_COUNTER_TX        : in std_logic_vector(2 downto 0);
   NACK_COUNTER_TX       : in std_logic_vector(2 downto 0);
   FCT_COUNTER_TX        : in std_logic_vector(3 downto 0);
   ACK_COUNTER_RX        : in std_logic_vector(2 downto 0);
   NACK_COUNTER_RX       : in std_logic_vector(2 downto 0);
   FCT_COUNTER_RX        : in std_logic_vector(3 downto 0);
   FULL_COUNTER_RX       : in std_logic_vector(1 downto 0);
   RETRY_COUNTER_RX      : in std_logic_vector(1 downto 0);
   CURRENT_TIME_SLOT     : in std_logic_vector(7 downto 0);
   LINK_RST_ASSERTED     : in std_logic;                                         -- Link has been reseted
   ACK_SEQ_NUM           : in std_logic_vector(7 downto 0);
   NACK_SEQ_NUM          : in std_logic_vector(7 downto 0);

   -- from the LANE
   LANE_STATE            : in std_logic_vector(C_LANESTATE_WIDTH-1 downto 0);    -- Lane state field
   RX_ERROR_CNT          : in std_logic_vector(C_RX_ERR_CNT_WIDTH-1 downto 0);   -- RX Error Counter
   RX_ERROR_OVF          : in std_logic;                                         -- RX Error Overflow
   LOSS_SIGNAL           : in std_logic;                                         -- Far-end lost Signal
   FAR_END_CAPA          : in std_logic_vector(C_FAR_CAPA_WIDTH-1 downto 0);     -- Far-end Capablities
   RX_POLARITY           : in std_logic;                                         -- RX Polarity

   -- to the DUT
   RST_DUT_N             : out std_logic;                                         -- Reset DUT (active low)
   DL_EN                 : out std_logic;                                         -- Lane injector enable command
   LANE_SPY_EN           : out std_logic;                                         -- Lane spy enable command

   -- from the DUT
   RESET_PARAM_DL        : in std_logic                                           -- Reset configuration parameters control
   );
end DATA_LINK_CONFIGURATOR;

------------------------------------------------------------------------------------------------------------------
--                                                  ARCHITECTURE                                                --
------------------------------------------------------------------------------------------------------------------
architecture rtl of DATA_LINK_CONFIGURATOR is
---------------------------------------
-- TYPES
---------------------------------------
   type axi_wr_state_t is (IDLE_WAIT_WR_ADDR, WR_RESPONSE);                           -- Write states for FSM declaration
   type axi_rd_state_t is (IDLE_WAIT_RD_ADDR, RD_RESPONSE);                           -- Read states for FSM declaration

---------------------------------------
-- SIGNAL DECLARATION
---------------------------------------
   signal axi_wr_state : axi_wr_state_t;
   signal axi_rd_state : axi_rd_state_t;
   -- Registers
   ------------
   signal reg_dl_param     : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link parameters register
   signal reg_dl_err_mngt  : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link error management register
   signal reg_dl_status_1  : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link status register
   signal reg_dl_status_2  : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link status register
   signal reg_dl_qos_1     : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link status register
   signal reg_dl_qos_2     : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Data Link status register
   signal reg_lane_param   : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Lane parameters register
   signal reg_lane_status  : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Lane status register
   signal reg_phy_param    : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- PHY parameters register
   signal reg_global       : std_logic_vector(G_DATA_WIDTH-1 downto 0);               -- Global register
   -- internal signals dl
   ------------
   signal vc_credit_i           :  std_logic_vector(G_CHANNEL_NUMBER-1 downto 0);     -- Up if each corresponding virtual channel has credit in the far-end input buffer
   signal fct_credit_overflow_i :  std_logic_vector(G_CHANNEL_NUMBER-1 downto 0);     -- Up if each corresponding virtual channel credit counter overflowed
   signal crc_long_error_i      :  std_logic;                                         -- RX error in CRC-16bit
   signal crc_short_error_i     :  std_logic;                                         -- RX error in CRC-8bit
   signal frame_error_i        :  std_logic;                                          -- RX frame error
   signal seq_error_i           :  std_logic;                                         -- RX SEQUENCE_NUMBER error
   signal far_end_link_rst_i    :  std_logic;                                         -- Far-end Link reset status
   signal seq_number_tx_i       :  std_logic_vector(7 downto 0);                      -- SEQ_NUMBER in transmission
   signal seq_number_rx_i       :  std_logic_vector(7 downto 0);                      -- SEQ_NUMBER in reception
   signal input_buffer_ovfl_i   :  std_logic_vector(7 downto 0);                      -- Up if each corresponding virtual channel input buffer overflowed
   -- internal signals lane and phy
   ------------
   signal lane_start_pulse : std_logic;                                               -- SpaceFibre lane start initialization signal pulsed

   signal lane_state_i     : std_logic_vector(C_LANESTATE_WIDTH-1 downto 0);          -- Lane state field
   signal rx_error_cnt_i   : std_logic_vector(C_RX_ERR_CNT_WIDTH-1 downto 0);         -- RX Error Counter
   signal rx_error_ovf_i   : std_logic;                                               -- RX Error Overflow
   signal loss_signal_i    : std_logic;                                               -- Far-end lost Signal
   signal far_end_capa_i   : std_logic_vector(C_FAR_CAPA_WIDTH-1 downto 0);           -- Far-end Capablities
   signal rx_polarity_i    : std_logic;                                               -- RX Polarity
   -- inputs resynchronization
   signal outputs_to_sync_lane  : std_logic_vector(13 downto 0);                      -- Signal to Lane layer of the DUT before synchronization
   signal outputs_to_dut_lane   : std_logic_vector(13 downto 0);                      -- Signal to Lane layer of the DUT after synchronization

   signal outputs_to_sync_dl  : std_logic_vector(22 downto 0);                        -- Signal to Data Link layer of the DUT before synchronization
   signal outputs_to_dut_dl   : std_logic_vector(22 downto 0);                        -- Signal to Data Link layer of the DUT after synchronization
   -- inputs resynchronization
   signal inputs_to_sync   : std_logic_vector(149 downto 0);                          -- Signal from the DUT before synchronization
   signal inputs_to_model  : std_logic_vector(149 downto 0);                          -- Signal from the DUT after synchronization

   signal frame_tx_i           : std_logic_vector(8 downto 0);                        -- Frame Tx 
   signal frame_finished_i     : std_logic_vector(8 downto 0);                        -- Frame Finished
   signal data_cnt_tx_i        : std_logic_vector(6 downto 0);                        -- Data Cnt TX
   signal data_cnt_rx_i        : std_logic_vector(6 downto 0);                        -- Data Cnt RX
   signal ack_counter_tx_i     : std_logic_vector(2 downto 0);                        -- Ack Counter TX
   signal nack_counter_tx_i    : std_logic_vector(2 downto 0);                        -- Nack Counter TX
   signal fct_counter_tx_i     : std_logic_vector(3 downto 0);                        -- Fct Counter TX
   signal ack_counter_rx_i     : std_logic_vector(2 downto 0);                        -- Ack Counter RX
   signal nack_counter_rx_i    : std_logic_vector(2 downto 0);                        -- Nack Counter RX
   signal fct_counter_rx_i     : std_logic_vector(3 downto 0);                        -- Fct Counter RX
   signal full_counter_rx_i    : std_logic_vector(1 downto 0);                        -- Full Counter RX
   signal retry_counter_rx_i   : std_logic_vector(1 downto 0);                        -- Retry Counter RX
   signal current_time_slot_i  : std_logic_vector(7 downto 0);                        -- Current Time-Slot
   signal link_rst_asserted_i  : std_logic;                                           -- Link Rst Asserted
   signal reset_param_dl_i     : std_logic;                                           -- Reset Param DL
   signal clear_error_flag     : std_logic;                                           -- Clear Error Flag
   signal ack_seq_num_i        : std_logic_vector(7 downto 0);                        -- Ack Seq num
   signal nack_seq_num_i       : std_logic_vector(7 downto 0);                        -- Nack Seq num
   signal dl_en_i              : std_logic;                                           -- Injector enable
   signal lane_spy_en_i        : std_logic;                                           -- Lane Spy enable

   begin
---------------------------------------
-- SIGNAL CONNECTION
---------------------------------------

    -- Parameter from Configurator to Lane
    outputs_to_sync_lane(0)           <= reg_lane_param(C_LANESTART_BTFD) or lane_start_pulse;
    outputs_to_sync_lane(1)           <= reg_lane_param(C_AUTOSTART_BTFD);
    outputs_to_sync_lane(2)           <= reg_lane_param(C_LANERESET_BTFD);
    outputs_to_sync_lane(3)           <= reg_lane_param(C_PARALLEL_LPB_BTFD);
    outputs_to_sync_lane(11 downto 4) <= reg_lane_param(C_STDBREASON_MAX_BTFD downto C_PARALLEL_LPB_BTFD +1);

    LANE_START                   <= outputs_to_dut_lane(0);
    AUTOSTART                    <= outputs_to_dut_lane(1);
    LANE_RESET                   <= outputs_to_dut_lane(2);
    PARALLEL_LOOPBACK_EN         <= outputs_to_dut_lane(3);
    STANDBY_REASON               <= outputs_to_dut_lane(11 downto 4);

    -- Parameter from Configurator to Phy
    outputs_to_sync_lane(13)          <= reg_phy_param(C_FAR_END_LPB_BTFD);
    outputs_to_sync_lane(12)          <= reg_phy_param(C_NEAR_END_LPB_BTFD);

    NEAR_END_SERIAL_LB_EN        <= outputs_to_dut_lane(12);
    FAR_END_SERIAL_LB_EN         <= outputs_to_dut_lane(13);

    -- Parameter from Configurator to Data Link
    outputs_to_sync_dl(0)           <= reg_dl_param(C_INTERFACE_RST_BTFD);
    outputs_to_sync_dl(1)           <= reg_dl_param(C_LINK_RST_BTFD);
    outputs_to_sync_dl(2)           <= reg_dl_param(C_NACK_RST_EN_BTFD);
    outputs_to_sync_dl(3)           <= reg_dl_param(C_NACK_RST_MODE_BTFD);
    outputs_to_sync_dl(12 downto 4) <= reg_dl_param(C_PAUSE_VC_BTFD downto C_NACK_RST_MODE_BTFD + 1);
    outputs_to_sync_dl(20 downto 13) <= reg_dl_param(C_CONTINUOUS_VC_BTFD downto C_PAUSE_VC_BTFD + 1);

    outputs_to_sync_dl(21)            <= dl_en_i;
    outputs_to_sync_dl(22)            <= lane_spy_en_i;
    clear_error_flag              <= reg_dl_param (C_CLEAR_ERROR_FLAG_BTFD);

    INTERFACE_RST                <= outputs_to_dut_dl(0);
    LINK_RST                     <= outputs_to_dut_dl(1);
    NACK_RST_EN                  <= outputs_to_dut_dl(2);
    NACK_RST_MODE                <= outputs_to_dut_dl(3);
    PAUSE_VC                     <= outputs_to_dut_dl(12 downto 4);
    CONTINUOUS_VC                <= outputs_to_dut_dl(20 downto 13);

    DL_EN                        <= outputs_to_dut_dl(21);
    LANE_SPY_EN                  <= outputs_to_dut_dl(22);

    -- Status from Lane  to Configurator
    inputs_to_sync(3 downto 0)              <= LANE_STATE;
    inputs_to_sync(11 downto 4)             <= RX_ERROR_CNT;
    inputs_to_sync(12)                      <= RX_ERROR_OVF;
    inputs_to_sync(13)                      <= LOSS_SIGNAL;
    inputs_to_sync(21 downto 14)            <= FAR_END_CAPA;
    inputs_to_sync(22)                      <= RX_POLARITY;

    lane_state_i                 <= inputs_to_model(3 downto 0);
    rx_error_cnt_i               <= inputs_to_model(11 downto 4);
    rx_error_ovf_i               <= inputs_to_model(12);
    loss_signal_i                <= inputs_to_model(13);
    far_end_capa_i               <= inputs_to_model(21 downto 14);
    rx_polarity_i                <= inputs_to_model(22);


   -- Status and QoS from Data Link to Configurator
    inputs_to_sync(30 downto 23)                 <= VC_CREDIT;
    inputs_to_sync(38 downto 31)                 <= FCT_CREDIT_OVERFLOW;
    inputs_to_sync(39)                           <= CRC_LONG_ERROR;
    inputs_to_sync(40)                           <= CRC_SHORT_ERROR;
    inputs_to_sync(41)                           <= FRAME_ERROR;
    inputs_to_sync(42)                           <= SEQ_ERROR;
    inputs_to_sync(43)                           <= FAR_END_LINK_RST;
    inputs_to_sync(51 downto 44)                 <= SEQ_NUMBER_TX;
    inputs_to_sync(59 downto 52)                 <= SEQ_NUMBER_RX;
    inputs_to_sync(67 downto 60)                 <= INPUT_BUFFER_OVFL;
    inputs_to_sync(76 downto 68)                 <= FRAME_TX;
    inputs_to_sync(85 downto 77)                 <= FRAME_FINISHED;
    inputs_to_sync(92 downto 86)                 <= DATA_CNT_TX;
    inputs_to_sync(99 downto 93)                 <= DATA_CNT_RX;
    inputs_to_sync(102 downto 100)               <= ACK_COUNTER_TX;
    inputs_to_sync(105 downto 103)               <= NACK_COUNTER_TX;
    inputs_to_sync(109 downto 106)               <= FCT_COUNTER_TX;
    inputs_to_sync(112 downto 110)               <= ACK_COUNTER_RX;
    inputs_to_sync(115 downto 113)               <= NACK_COUNTER_RX;
    inputs_to_sync(119 downto 116)               <= FCT_COUNTER_RX;
    inputs_to_sync(121 downto 120)               <= FULL_COUNTER_RX;
    inputs_to_sync(123 downto 122)               <= RETRY_COUNTER_RX;
    inputs_to_sync(131 downto 124)               <= CURRENT_TIME_SLOT;
    inputs_to_sync(132)                          <= LINK_RST_ASSERTED;
    inputs_to_sync(140 downto 133)               <= ACK_SEQ_NUM;
    inputs_to_sync(148 downto 141)               <= NACK_SEQ_NUM;

    vc_credit_i                 <= inputs_to_model(30 downto 23);
    fct_credit_overflow_i       <= inputs_to_model(38 downto 31);
    crc_long_error_i            <= inputs_to_model(39);
    crc_short_error_i           <= inputs_to_model(40);
    frame_error_i               <= inputs_to_model(41);
    seq_error_i                 <= inputs_to_model(42);
    far_end_link_rst_i          <= inputs_to_model(44);
    seq_number_tx_i             <= inputs_to_model(51 downto 44);
    seq_number_rx_i             <= inputs_to_model(59 downto 52);
    input_buffer_ovfl_i         <= inputs_to_model(67 downto 60) or reg_dl_status_2(C_INPUT_BUFFER_OVERFLW_BTFD downto C_FAR_END_LINK_RST_BTFD + 1);
    frame_tx_i                  <= inputs_to_model(76 downto 68);
    frame_finished_i            <= inputs_to_model(85 downto 77);
    data_cnt_tx_i               <= inputs_to_model(92 downto 86);
    data_cnt_rx_i               <= inputs_to_model(99 downto 93);
    ack_counter_tx_i            <= inputs_to_model(102 downto 100);
    nack_counter_tx_i           <= inputs_to_model(105 downto 103);
    fct_counter_tx_i            <= inputs_to_model(109 downto 106);
    ack_counter_rx_i            <= inputs_to_model(112 downto 110);
    nack_counter_rx_i           <= inputs_to_model(115 downto 113);
    fct_counter_rx_i            <= inputs_to_model(119 downto 116);
    full_counter_rx_i           <= inputs_to_model(121 downto 120);
    retry_counter_rx_i          <= inputs_to_model(123 downto 122);
    current_time_slot_i         <= inputs_to_model(131 downto 124);
    link_rst_asserted_i         <= inputs_to_model(132);
    ack_seq_num_i               <= inputs_to_model(140 downto 133);
    nack_seq_num_i              <= inputs_to_model(148 downto 141);

    -- Parameters reset from Data Link to configurator
    inputs_to_sync(149)         <= RESET_PARAM_DL;
    reset_param_dl_i            <= inputs_to_model(149);

   lane_start_pulse             <= reg_lane_param(C_LANESTART_PULSE_BTFD);
   RST_DUT_N                    <= reg_global(C_RST_DUT_BTFD);
   dl_en_i                      <= reg_global(C_DL_EN_BTFD);
   lane_spy_en_i                <= reg_global(C_LANE_SPY_EN_BTFD);

---------------------------------------
-- INSTANCIATION
---------------------------------------
  ---------------------------------------------------------------------------
  -- INSTANCE: I_RESYNC_OUT_LANE
  -- Description : Resynchronize signals from the model at CLK to the CLK_TX clock
  ---------------------------------------------------------------------------
  I_RESYNC_OUT_LANE: entity work.resync_double
  generic map (
   VECTOR_SIZE => outputs_to_sync_lane'length
  )
  port map (
   -- system signals
   clk    => CLK_TX,                                                               --- main clock
   rst_n  => RST_TXCLK_N,                                                          --- main reset (active low)
   -- I/Os
   input  => outputs_to_sync_lane,                                                 --- vector to synchronize
   output => outputs_to_dut_lane                                                   --- double synchronized vector
  );
  ---------------------------------------------------------------------------
  -- INSTANCE: I_RESYNC_OUT_DL
  -- Description : Resynchronize signals from the model at CLK to the CLK_TX clock
  ---------------------------------------------------------------------------
  I_RESYNC_OUT_DL: entity work.resync_double
  generic map (
   VECTOR_SIZE => outputs_to_sync_dl'length
  )
  port map (
   -- system signals
   clk    => CLK_DL,                                                               --- main clock
   rst_n  => RST_N_DL,                                                             --- main reset (active low)
   -- I/Os
   input  => outputs_to_sync_dl,                                                   --- vector to synchronize
   output => outputs_to_dut_dl                                                     --- double synchronized vector
  );
  ---------------------------------------------------------------------------
  -- INSTANCE: I_RESYNC_IN
  -- Description : Resynchronize signals from the DUT at CLK_TX to the CLK clock
   ---------------------------------------------------------------------------
  I_RESYNC_IN: entity work.resync_double
  generic map (
   VECTOR_SIZE => inputs_to_sync'length
  )
  port map (
   -- system signals
   clk    => CLK,                                                                  --- main clock
   rst_n  => RST_N,                                                                --- main reset (active low)
   -- I/Os
   input  => inputs_to_sync,                                                       --- vector to synchronize
   output => inputs_to_model                                                       --- double synchronized vector
  );
---------------------------------------
-- PROCESS
---------------------------------------
   ---------------------------------------------------------------------------
   -- PROCESS: P_AXI_READ
   -- Description : AXI4 Lite reading process
   ---------------------------------------------------------------------------
   P_AXI_READ : process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N ='0') then
         axi_rd_state    <= IDLE_WAIT_RD_ADDR;
         S_AXI_ARREADY   <= '1';               -- Ready for new request
         S_AXI_RRESP     <= "00";              -- OKAY default response
         S_AXI_RDATA     <= (others => '0');   -- Default data at zero
         S_AXI_RVALID    <= '0';               -- Default read validity at zero
      elsif rising_edge(CLK) then
         case axi_rd_state is
            -- Waiting for a read request
            when IDLE_WAIT_RD_ADDR =>
               S_AXI_ARREADY <= '1';     -- Ready for new read request
               if (S_AXI_ARVALID = '1') then
                   S_AXI_ARREADY <= '0'; -- Ready signal deasserted to indicate request processing
                   -- Parameters lane register address
                   if (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_LANE_PARAM) then
                       S_AXI_RDATA  <= reg_lane_param;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Status lane register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_LANE_STATUS) then
                       S_AXI_RDATA  <= reg_lane_status;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Parameters PHY register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_PHY_PARAM) then
                       S_AXI_RDATA  <= reg_phy_param;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Parameters DL register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_PARAM) then
                       S_AXI_RDATA  <= reg_dl_param;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Status DL register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_STATUS_1) then
                      S_AXI_RDATA  <= reg_dl_status_1;
                      S_AXI_RRESP  <= "00";
                      S_AXI_RVALID <= '1';
                      axi_rd_state <= RD_RESPONSE;
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_STATUS_2) then
                      S_AXI_RDATA  <= reg_dl_status_2;
                      S_AXI_RRESP  <= "00";
                      S_AXI_RVALID <= '1';
                      axi_rd_state <= RD_RESPONSE;
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_QOS_1) then
                      S_AXI_RDATA  <= reg_dl_qos_1;
                      S_AXI_RRESP  <= "00";
                      S_AXI_RVALID <= '1';
                      axi_rd_state <= RD_RESPONSE;
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_QOS_2) then
                      S_AXI_RDATA  <= reg_dl_qos_2;
                      S_AXI_RRESP  <= "00";
                      S_AXI_RVALID <= '1';
                      axi_rd_state <= RD_RESPONSE;
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_ERR_MNGT) then
                        S_AXI_RDATA  <= reg_dl_err_mngt;
                        S_AXI_RRESP  <= "00";
                        S_AXI_RVALID <= '1';
                        axi_rd_state <= RD_RESPONSE;
                   -- Global register address
                   elsif (S_AXI_ARADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_GLOBAL) then
                       S_AXI_RDATA  <= reg_global;
                       S_AXI_RRESP  <= "00";
                       S_AXI_RVALID <= '1';
                       axi_rd_state <= RD_RESPONSE;
                   -- Unrecognized address
                   else
                       S_AXI_RDATA  <= (others => '0');   -- Default response data
                       S_AXI_RRESP  <= "10";              -- Error response (SLVERR)
                       S_AXI_RVALID <= '1';               -- Response valid
                       axi_rd_state <= RD_RESPONSE;       -- Send the error response
                   end if;
               -- No read request received
               else
                   axi_rd_state <= IDLE_WAIT_RD_ADDR;
               end if;
            -- Responding to the read request
            when RD_RESPONSE =>
               -- Waiting for data reception confirmation from the master
               if (S_AXI_RREADY = '1') then
                   S_AXI_RVALID  <= '0';               -- Deassertion of response validity
                   S_AXI_RDATA   <= (others => '0');   -- Data reset
                   S_AXI_RRESP   <= "00";              -- Default OKAY response
                   axi_rd_state <= IDLE_WAIT_RD_ADDR;
               -- Wait until the master's reception confirmation is received
               else
                   axi_rd_state <= RD_RESPONSE;
               end if;
            -- Unrecognized state, return to IDLE state
            when others =>
               axi_rd_state <= IDLE_WAIT_RD_ADDR;
         end case;
      end if;
   end process P_AXI_READ;
   ---------------------------------------------------------------------------
   -- PROCESS: P_AXI_WRITE
   -- Description : AXI4 Lite writing process
   ---------------------------------------------------------------------------
   P_AXI_WRITE: process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N = '0' ) then
         axi_wr_state    <= IDLE_WAIT_WR_ADDR;
         S_AXI_AWREADY   <= '1';                 -- Ready for new request
         S_AXI_WREADY    <= '1';                 -- Ready to receive write data
         S_AXI_BRESP     <= "00";                -- OKAY default response
         S_AXI_BVALID    <= '0';                 -- Default write response validity
         reg_dl_param    <= init_dl_dl_param;
         reg_lane_param  <= init_lc_lane_param;
         reg_phy_param   <= init_lc_phy_param;
         reg_global      <= init_lc_global;
      elsif rising_edge(CLK) then
         if (lane_start_pulse ='1') then
            reg_lane_param(C_LANESTART_PULSE_BTFD)  <= '0';  -- Reset model start bit
         end if;
         if (reset_param_dl_i = '1') then                    -- Configuration reset from data link
            reg_dl_param                            <= init_dl_dl_param;
            reg_lane_param                          <= init_lc_lane_param;
            reg_phy_param                           <= init_lc_phy_param;
         end if;
         if link_rst_asserted_i = '1' then                   -- Link reset command from data link
            reg_dl_param(C_LINK_RST_ASSERTED_BTFD)  <= link_rst_asserted_i;
         end if;
         if clear_error_flag = '1' then                      -- Flag to clear the error counter
            reg_dl_param(C_CLEAR_ERROR_FLAG_BTFD)   <= '0';
         end if;
         case axi_wr_state is
            -- Waiting for a write request
            when IDLE_WAIT_WR_ADDR =>
               S_AXI_AWREADY    <= '1';              -- Ready for new request
               S_AXI_WREADY     <= '1';
               if (S_AXI_AWVALID = '1' and S_AXI_WVALID ='1') then
                  S_AXI_AWREADY   <= '0';           -- Ready signals deasserted to indicate request processing
                  S_AXI_WREADY    <= '0';
                  -- Parameters lane register address
                  if (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_LANE_PARAM) then
                     reg_lane_param <= S_AXI_WDATA; -- Write lane parameters
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Parameters phy register address
                  elsif (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_PHY_PARAM) then
                     reg_phy_param  <= S_AXI_WDATA; -- Write phy parameters
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Parameter DL register address
                  elsif (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_DL_PARAM) then
                     reg_dl_param   <= S_AXI_WDATA; -- Write DL parameters
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Global control register address
                  elsif (S_AXI_AWADDR(C_SLAVE_ADDR_WIDTH-1 downto 0) = C_ADDR_DL_GLOBAL) then
                     reg_global     <= S_AXI_WDATA; -- Write global signals
                     S_AXI_BRESP    <= "00";        -- OKAY response
                     S_AXI_BVALID   <= '1';         -- Valid response
                     axi_wr_state   <= WR_RESPONSE;
                  -- Unrecognized address
                  else
                     S_AXI_BRESP  <= "10";          -- Error response (SLVERR)
                     S_AXI_BVALID <= '1';           -- Response valid
                     axi_wr_state <= WR_RESPONSE;
                  end if;
               -- No write request received
               else
                  axi_wr_state <= IDLE_WAIT_WR_ADDR;
               end if;
            -- Responding to the write request
            when WR_RESPONSE =>
               -- Waiting for response reception confirmation from the master
               if (S_AXI_BREADY  = '1') then
                  S_AXI_BVALID    <= '0';           -- Reset response validity
                  S_AXI_BRESP     <= "00";          -- Default OKAY response
                  axi_wr_state <= IDLE_WAIT_WR_ADDR;
               -- Wait until the master's reception confirmation is received
               else
                  axi_wr_state <= WR_RESPONSE;
               end if;
            -- Unrecognized state, return to IDLE state
            when others =>
                axi_wr_state <= IDLE_WAIT_WR_ADDR;
         end case;
      end if;
   end process P_AXI_WRITE;
   ---------------------------------------------------------------------------
   -- PROCESS: P_STATUS
   -- Description : update status register
   ---------------------------------------------------------------------------
   P_STATUS : process(CLK, RST_N)
   begin
      -- Reset
      if (RST_N ='0') then
         reg_lane_status                                                                  <= (others => '0');
         reg_dl_status_1                                                                  <= (others => '0');
         reg_dl_status_2                                                                  <= (others => '0');
         reg_dl_err_mngt                                                                  <= (others => '0');
      elsif rising_edge(CLK) then
         reg_lane_status(C_RX_POLARITY_BTFD)                                              <= rx_polarity_i;
         reg_lane_status(C_FAR_CAPA_MAX_BTFD downto C_FAR_LOST_SIG_BTFD+1)                <= far_end_capa_i;
         reg_lane_status(C_FAR_LOST_SIG_BTFD)                                             <= loss_signal_i;
         reg_lane_status(C_RX_ERR_OVF_BTFD)                                               <= rx_error_ovf_i;
         reg_lane_status(C_RX_ERR_CNT_MAX_BTFD downto C_LANESTATE_MAX_BTFD+1)             <= rx_error_cnt_i;
         reg_lane_status(C_LANESTATE_MAX_BTFD downto 0)                                   <= lane_state_i;
         reg_dl_status_1(C_SEQ_NUMBER_TX_BTFD downto 0)                                   <= seq_number_tx_i;
         reg_dl_status_1(C_SEQ_NUMBER_RX_BTFD downto C_SEQ_NUMBER_TX_BTFD + 1)            <= seq_number_rx_i;
         reg_dl_status_1(C_VC_CREDIT_BTFD downto C_SEQ_NUMBER_RX_BTFD + 1)                <= vc_credit_i;
         reg_dl_status_1(C_FCT_CREDIT_OVERFLOW_BTFD downto C_VC_CREDIT_BTFD + 1)          <= fct_credit_overflow_i;
         if crc_long_error_i ='1' then    -- Stay up to be readable by the AXI interface, need tobe cleared manually
            reg_dl_status_2(C_CRC_LONG_ERROR_BTFD)                                        <= crc_long_error_i;
         end if;
         if crc_short_error_i = '1' then  -- Stay up to be readable by the AXI interface, need tobe cleared manually
            reg_dl_status_2(C_CRC_SHORT_ERROR_BTFD)                                       <= crc_short_error_i;
         end if;
         if frame_error_i = '1' then      -- Stay up to be readable by the AXI interface, need tobe cleared manually
            reg_dl_status_2(C_FRAME_ERROR_BTFD)                                           <= frame_error_i;
         end if;
         if seq_error_i = '1' then        -- Stay up to be readable by the AXI interface, need tobe cleared manually
            reg_dl_status_2(C_SEQ_ERROR_BTFD)                                             <= seq_error_i;
         end if;
         reg_dl_status_2(C_FAR_END_LINK_RST_BTFD)                                         <= far_end_link_rst_i;
         reg_dl_status_2(C_INPUT_BUFFER_OVERFLW_BTFD downto C_FAR_END_LINK_RST_BTFD + 1)  <= input_buffer_ovfl_i;
         reg_dl_qos_1(C_FRAME_FINISHED_BTFD downto 0)                                     <= frame_finished_i;
         reg_dl_qos_1(C_FRAME_TX_BTFD downto C_FRAME_FINISHED_BTFD + 1)                   <= frame_tx_i;
         reg_dl_qos_1(C_DATA_CNT_TX_BTFD downto C_FRAME_TX_BTFD + 1)                      <= data_cnt_tx_i;
         reg_dl_qos_1(C_DATA_CNT_RX_BTFD downto C_DATA_CNT_TX_BTFD + 1)                   <= data_cnt_rx_i;
         reg_dl_qos_2(C_ACK_COUNTER_TX_BTFD downto 0)                                     <= ack_counter_tx_i;
         reg_dl_qos_2(C_NACK_COUNTER_TX_BTFD downto C_ACK_COUNTER_TX_BTFD +1)             <= nack_counter_tx_i;
         reg_dl_qos_2(C_FCT_COUNTER_TX_BTFD downto C_NACK_COUNTER_TX_BTFD +1)             <= fct_counter_tx_i;
         reg_dl_qos_2(C_ACK_COUNTER_RX_BTFD downto C_FCT_COUNTER_TX_BTFD +1)              <= ack_counter_rx_i;
         reg_dl_qos_2(C_NACK_COUNTER_RX_BTFD downto C_ACK_COUNTER_RX_BTFD +1)             <= nack_counter_rx_i;
         reg_dl_qos_2(C_FCT_COUNTER_RX_BTFD downto C_NACK_COUNTER_RX_BTFD +1)             <= fct_counter_rx_i;
         reg_dl_qos_2(C_FULL_COUNTER_RX_BTFD downto C_FCT_COUNTER_RX_BTFD + 1)            <= full_counter_rx_i;
         reg_dl_qos_2(C_RETRY_COUNTER_RX_BTFD downto C_FULL_COUNTER_RX_BTFD + 1)          <= retry_counter_rx_i;
         reg_dl_qos_2(C_CURRENT_TIME_SLOT_BTFD downto C_RETRY_COUNTER_RX_BTFD + 1)        <= current_time_slot_i;
         reg_dl_err_mngt(C_ACK_SEQ_NUM_BTFD downto 0)                                     <= ack_seq_num_i;
         reg_dl_err_mngt(C_NACK_SEQ_NUM_BTFD downto C_ACK_SEQ_NUM_BTFD + 1)               <= nack_seq_num_i;
         if clear_error_flag = '1' then  -- Manual clear of error counter with clear_error_flag
            reg_dl_status_2(C_CRC_LONG_ERROR_BTFD)                                           <= '0';
            reg_dl_status_2(C_CRC_SHORT_ERROR_BTFD)                                          <= '0';
            reg_dl_status_2(C_FRAME_ERROR_BTFD)                                              <= '0';
            reg_dl_status_2(C_SEQ_ERROR_BTFD)                                                <= '0';
            reg_dl_status_2(C_INPUT_BUFFER_OVERFLW_BTFD downto C_FAR_END_LINK_RST_BTFD + 1)  <= (others => '0');
         end if;
      end if;
   end process P_STATUS;
end rtl;
