-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 18/06/2025
--
-- Description : This module allows realigning the beginnings of words so
--               that they start on byte 0 or 4.
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
  use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_word_alignment is
  port (
    RST_N                   : in  std_logic;                                   --! Global reset. Active low
    CLK                     : in  std_logic;                                   --! Clock generated by HSSL IP
    -- ppl_64_rx_sync_fsm (PLRSF) interface
    DATA_RX_PLWA            : out std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data to lane_ctrl_word_detect
    VALID_K_CHARAC_PLWA     : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags to lane_ctrl_word_detect
    DATA_RDY_PLWA           : out std_logic;                                   --! Data valid flag to lane_ctrl_word_detect
    INVALID_CHAR_PLWA       : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Invalid character flags from PLWA
    DISPARITY_ERR_PLWA      : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Disparity error flags from PLWA
    RX_WORD_IS_ALIGNED_PLWA : out std_logic;                                   --! RX word is aligned from PLWA
    COMMA_DET_PLWA          : out std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flag indicates that a comma is detected on the word receive from PLWA
    LOSS_OF_SIGNAL_PLWA     : out  std_logic;                                  --! Loss of signal flag from PLWA
    -- HSSL IP interface
    DATA_RX_HSSL            : in  std_logic_vector(C_DATA_WIDTH-1 downto 0);   --! 64-bit data from HSSL IP
    VALID_K_CHARAC_HSSL     : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! 8-bit valid K character flags from HSSL IP
    INVALID_CHAR_HSSL       : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Invalid character flags from HSSL IP
    DISPARITY_ERR_HSSL      : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Disparity error flags from HSSL IP
    RX_WORD_IS_ALIGNED_HSSL : in  std_logic;                                   --! RX word is aligned from HSSL IP
    RX_VALID_REALIGN_HSSL : in  std_logic;                                   --! RX word is aligned from HSSL IP
    COMMA_DET_HSSL          : in  std_logic_vector(C_K_CHAR_WIDTH-1 downto 0); --! Flag indicates that a comma is detected on the word receive
    LOSS_OF_SIGNAL_HSSL     : in  std_logic                                   --! Loss of signal flag from HSSL IP
  );
end ppl_64_word_alignment;

architecture rtl of ppl_64_word_alignment is
---------------------------------------------------------
----- Type declaration -----
---------------------------------------------------------
type rx_word_align_fsm_type is (
   INIT_ST,  --! INIT state of the FSM waiting for alignment
   WAITING_COMMA_ST,
   ALIGNED_ST --! Checking data to validate synchronization state
   );
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
  signal current_state               : rx_word_align_fsm_type;
  signal reg_data                    : std_logic_vector(C_DATA_WIDTH-1 downto 0);
  signal reg_k_char                  : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal reg_invalid_k_char          : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal reg_disp_err                : std_logic_vector(C_K_CHAR_WIDTH-1 downto 0);
  signal alignment_byte              : unsigned(C_K_CHAR_WIDTH-1 downto 0);
begin
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_rx_realignment
--! Aligns the words so that they are at the beginning of the bus.
---------------------------------------------------------
  p_rx_realignment: process(CLK,RST_N)
  begin
    if RST_N = '0' then
      DATA_RX_PLWA        <= (others => '0');
      VALID_K_CHARAC_PLWA <= (others => '0');
      DATA_RDY_PLWA       <= '0';
      INVALID_CHAR_PLWA   <= (others => '0');
      DISPARITY_ERR_PLWA  <= (others => '0');
      alignment_byte      <= (others => '0');
      reg_data            <= (others => '0');
      reg_k_char          <= (others => '0');
      reg_invalid_k_char  <= (others => '0');
      reg_disp_err        <= (others => '0');
      current_state       <= INIT_ST;
    elsif rising_edge(CLK) then
      case current_state is
        when INIT_ST  =>
          -- Word is aligned
          if RX_WORD_IS_ALIGNED_HSSL ='1' and RX_VALID_REALIGN_HSSL= '1' then
            current_state  <= WAITING_COMMA_ST;
          end if;

        when WAITING_COMMA_ST =>
          -- Word is aligned
          if RX_WORD_IS_ALIGNED_HSSL ='1' then
            -- Comma on byte 7
            if COMMA_DET_HSSL(7) = '1'  then
              alignment_byte      <= "10000000";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(7*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 7*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(7-1 downto 0) & reg_k_char(7);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(7-1 downto 0) & reg_invalid_k_char(7);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(7-1 downto 0) & reg_disp_err(7);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 6
            elsif COMMA_DET_HSSL(6) = '1'  then
              alignment_byte      <= "01000000";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(6*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 6*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(6-1 downto 0) & reg_k_char(7 downto 6);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(6-1 downto 0) & reg_invalid_k_char(7 downto 6);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(6-1 downto 0) & reg_disp_err(7 downto 6);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 5
            elsif COMMA_DET_HSSL(5) = '1' then
              alignment_byte      <= "00100000";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(5*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 5*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(5-1 downto 0) & reg_k_char(7 downto 5);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(5-1 downto 0) & reg_invalid_k_char(7 downto 5);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(5-1 downto 0) & reg_disp_err(7 downto 5);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 4
            elsif COMMA_DET_HSSL(4) = '1' then
              alignment_byte      <= "00010000";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(4*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 4*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(4-1 downto 0) & reg_k_char(7 downto 4);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(4-1 downto 0) & reg_invalid_k_char(7 downto 4);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(4-1 downto 0) & reg_disp_err(7 downto 4);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 3
            elsif COMMA_DET_HSSL(3) = '1' then
              alignment_byte      <= "00001000";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(3*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 3*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(3-1 downto 0) & reg_k_char(7 downto 3);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(3-1 downto 0) & reg_invalid_k_char(7 downto 3);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(3-1 downto 0) & reg_disp_err(7 downto 3);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 2
            elsif COMMA_DET_HSSL(2) = '1' then
              alignment_byte      <= "00000100";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(2*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 2*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(2-1 downto 0) & reg_k_char(7 downto 2);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(2-1 downto 0) & reg_invalid_k_char(7 downto 2);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(2-1 downto 0) & reg_disp_err(7 downto 2);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 1
            elsif COMMA_DET_HSSL(1) = '1' then
              alignment_byte      <= "00000010";
              reg_data            <= DATA_RX_HSSL;
              DATA_RX_PLWA        <= DATA_RX_HSSL(1*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 1*8);
              reg_k_char          <= VALID_K_CHARAC_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(1-1 downto 0) & reg_k_char(7 downto 1);
              reg_invalid_k_char  <= INVALID_CHAR_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL(1-1 downto 0) & reg_invalid_k_char(7 downto 1);
              reg_disp_err        <= DISPARITY_ERR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL(1-1 downto 0) & reg_disp_err(7 downto 1);
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- Comma on byte 0
            elsif COMMA_DET_HSSL(0) = '1' then
              alignment_byte      <= "00000001";
              DATA_RX_PLWA        <= DATA_RX_HSSL;
              VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL;
              INVALID_CHAR_PLWA   <= INVALID_CHAR_HSSL;
              DISPARITY_ERR_PLWA  <= DISPARITY_ERR_HSSL;
              DATA_RDY_PLWA       <= '1';
              current_state       <= ALIGNED_ST;
            -- No comma is detected
            else
              DATA_RX_PLWA        <= (others => '0');
              VALID_K_CHARAC_PLWA <= (others => '0');
              DATA_RDY_PLWA       <= '0';
              alignment_byte      <= (others => '0');
              reg_data            <= (others => '0');
              reg_k_char          <= (others => '0');
            end if;
          -- Word is not aligned
          else
            DATA_RX_PLWA        <= (others => '0');
            VALID_K_CHARAC_PLWA <= (others => '0');
            DATA_RDY_PLWA       <= '0';
            alignment_byte      <= (others => '0');
            reg_data            <= (others => '0');
            reg_k_char          <= (others => '0');
            current_state       <= INIT_ST;
          end if;

        when ALIGNED_ST  =>
          -- Word is aligned
          if RX_WORD_IS_ALIGNED_HSSL = '1' then
            -- When a comma is present, it is placed at the same position in the word
            if (std_logic_vector(alignment_byte(7 downto 4)) = COMMA_DET_HSSL(7 downto 4) or std_logic_vector(alignment_byte(3 downto 0)) = COMMA_DET_HSSL(7 downto 4))and
               (std_logic_vector(alignment_byte(7 downto 4)) = COMMA_DET_HSSL(3 downto 0) or std_logic_vector(alignment_byte(3 downto 0)) = COMMA_DET_HSSL(3 downto 0)) then
              -- Comma on byte 7
              if alignment_byte(7) = '1' then
                alignment_byte      <= "10000000";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(7*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 7*8)  ;
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(7-1 downto 0) & reg_k_char(7);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 6
              elsif alignment_byte(6) = '1' then
                alignment_byte      <= "01000000";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(6*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 6*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(6-1 downto 0) & reg_k_char(7 downto 6);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 5
              elsif alignment_byte(5) = '1' then
                alignment_byte      <= "00100000";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(5*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 5*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(5-1 downto 0) & reg_k_char(7 downto 5);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 4
              elsif alignment_byte(4) = '1' then
                alignment_byte      <= "00010000";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(4*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 4*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(4-1 downto 0) & reg_k_char(7 downto 4);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 3
              elsif alignment_byte(3) = '1' then
                alignment_byte      <= "00001000";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(3*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 3*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(3-1 downto 0) & reg_k_char(7 downto 3);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 2
              elsif alignment_byte(2) = '1' then
                alignment_byte      <= "00000100";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(2*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 2*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(2-1 downto 0) & reg_k_char(7 downto 2);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 1
              elsif alignment_byte(1) = '1' then
                alignment_byte      <= "00000010";
                reg_data            <= DATA_RX_HSSL;
                DATA_RX_PLWA        <= DATA_RX_HSSL(1*8-1 downto 0) & reg_data(C_K_CHAR_WIDTH*8-1 downto 1*8);
                reg_k_char          <= VALID_K_CHARAC_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL(1-1 downto 0) & reg_k_char(7 downto 1);
                DATA_RDY_PLWA       <= '1';
              -- Comma on byte 0
              elsif alignment_byte(0) = '1' then
                alignment_byte      <= "00000001";
                DATA_RX_PLWA        <= DATA_RX_HSSL;
                VALID_K_CHARAC_PLWA <= VALID_K_CHARAC_HSSL;
                DATA_RDY_PLWA       <= '1';
              else
                DATA_RX_PLWA        <= (others => '0');
                VALID_K_CHARAC_PLWA <= (others => '0');
                DATA_RDY_PLWA       <= '0';
                alignment_byte      <= (others => '0');
                reg_data            <= (others => '0');
                reg_k_char          <= (others => '0');
                current_state       <= WAITING_COMMA_ST;
              end if;
            -- Comma placed incorrectly
            else
              DATA_RX_PLWA        <= (others => '0');
              VALID_K_CHARAC_PLWA <= (others => '0');
              DATA_RDY_PLWA       <= '0';
              alignment_byte      <= (others => '0');
              reg_data            <= (others => '0');
              reg_k_char          <= (others => '0');
              current_state       <= WAITING_COMMA_ST;
            end if;
          -- Word is not aligned
          else
            DATA_RX_PLWA        <= (others => '0');
            VALID_K_CHARAC_PLWA <= (others => '0');
            DATA_RDY_PLWA       <= '0';
            alignment_byte      <= (others => '0');
            reg_data            <= (others => '0');
            reg_k_char          <= (others => '0');
            current_state       <= INIT_ST;
          end if;

        when others =>
          DATA_RX_PLWA        <= (others => '0');
          VALID_K_CHARAC_PLWA <= (others => '0');
          DATA_RDY_PLWA       <= '0';
          alignment_byte      <= (others => '0');
          reg_data            <= (others => '0');
          reg_k_char          <= (others => '0');
          current_state       <= INIT_ST;

        end case;
    end if;
  end process p_rx_realignment;
---------------------------------------------------------
-- Process: p_sync
--! Signals transfer
---------------------------------------------------------
  p_sync: process(CLK,RST_N)
  begin
    if RST_N = '0' then
      RX_WORD_IS_ALIGNED_PLWA <= '0';
      COMMA_DET_PLWA          <= (others => '0');
      LOSS_OF_SIGNAL_PLWA     <= '0';
    elsif rising_edge(CLK) then
      RX_WORD_IS_ALIGNED_PLWA <= RX_WORD_IS_ALIGNED_HSSL;
      COMMA_DET_PLWA          <= COMMA_DET_HSSL;
      LOSS_OF_SIGNAL_PLWA     <= LOSS_OF_SIGNAL_HSSL;
    end if;
  end process p_sync;

end architecture rtl;