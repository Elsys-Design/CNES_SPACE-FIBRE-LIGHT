// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC2_XBR2X4_DEFINES_VH
`else
`define B_NOC2_XBR2X4_DEFINES_VH

// Look-up table parameters
//

`define NOC2_XBR2X4_ADDR_N  119
`define NOC2_XBR2X4_ADDR_SZ 32
`define NOC2_XBR2X4_DATA_SZ 32

// Attribute addresses
//

`define NOC2_XBR2X4__REG_CLOCK_MUX    32'h00000000
`define NOC2_XBR2X4__REG_CLOCK_MUX_SZ 32

`define NOC2_XBR2X4__REG_HIGH_ID0_P_NMU    32'h00000001
`define NOC2_XBR2X4__REG_HIGH_ID0_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID10_P_NMU    32'h00000002
`define NOC2_XBR2X4__REG_HIGH_ID10_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID11_P_NMU    32'h00000003
`define NOC2_XBR2X4__REG_HIGH_ID11_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID12_P_NMU    32'h00000004
`define NOC2_XBR2X4__REG_HIGH_ID12_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID13_P_NMU    32'h00000005
`define NOC2_XBR2X4__REG_HIGH_ID13_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID14_P_NMU    32'h00000006
`define NOC2_XBR2X4__REG_HIGH_ID14_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID15_P_NMU    32'h00000007
`define NOC2_XBR2X4__REG_HIGH_ID15_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID16_P_NMU    32'h00000008
`define NOC2_XBR2X4__REG_HIGH_ID16_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID17_P_NMU    32'h00000009
`define NOC2_XBR2X4__REG_HIGH_ID17_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID18_P_NMU    32'h0000000a
`define NOC2_XBR2X4__REG_HIGH_ID18_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID19_P_NMU    32'h0000000b
`define NOC2_XBR2X4__REG_HIGH_ID19_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID1_P_NMU    32'h0000000c
`define NOC2_XBR2X4__REG_HIGH_ID1_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID20_P_NMU    32'h0000000d
`define NOC2_XBR2X4__REG_HIGH_ID20_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID21_P_NMU    32'h0000000e
`define NOC2_XBR2X4__REG_HIGH_ID21_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID22_P_NMU    32'h0000000f
`define NOC2_XBR2X4__REG_HIGH_ID22_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID23_P_NMU    32'h00000010
`define NOC2_XBR2X4__REG_HIGH_ID23_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID24_P_NMU    32'h00000011
`define NOC2_XBR2X4__REG_HIGH_ID24_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID25_P_NMU    32'h00000012
`define NOC2_XBR2X4__REG_HIGH_ID25_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID26_P_NMU    32'h00000013
`define NOC2_XBR2X4__REG_HIGH_ID26_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID27_P_NMU    32'h00000014
`define NOC2_XBR2X4__REG_HIGH_ID27_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID28_P_NMU    32'h00000015
`define NOC2_XBR2X4__REG_HIGH_ID28_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID29_P_NMU    32'h00000016
`define NOC2_XBR2X4__REG_HIGH_ID29_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID2_P_NMU    32'h00000017
`define NOC2_XBR2X4__REG_HIGH_ID2_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID30_P_NMU    32'h00000018
`define NOC2_XBR2X4__REG_HIGH_ID30_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID31_P_NMU    32'h00000019
`define NOC2_XBR2X4__REG_HIGH_ID31_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID32_P_NMU    32'h0000001a
`define NOC2_XBR2X4__REG_HIGH_ID32_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID33_P_NMU    32'h0000001b
`define NOC2_XBR2X4__REG_HIGH_ID33_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID34_P_NMU    32'h0000001c
`define NOC2_XBR2X4__REG_HIGH_ID34_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID35_P_NMU    32'h0000001d
`define NOC2_XBR2X4__REG_HIGH_ID35_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID36_P_NMU    32'h0000001e
`define NOC2_XBR2X4__REG_HIGH_ID36_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID37_P_NMU    32'h0000001f
`define NOC2_XBR2X4__REG_HIGH_ID37_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID38_P_NMU    32'h00000020
`define NOC2_XBR2X4__REG_HIGH_ID38_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID39_P_NMU    32'h00000021
`define NOC2_XBR2X4__REG_HIGH_ID39_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID3_P_NMU    32'h00000022
`define NOC2_XBR2X4__REG_HIGH_ID3_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID40_P_NMU    32'h00000023
`define NOC2_XBR2X4__REG_HIGH_ID40_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID41_P_NMU    32'h00000024
`define NOC2_XBR2X4__REG_HIGH_ID41_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID42_P_NMU    32'h00000025
`define NOC2_XBR2X4__REG_HIGH_ID42_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID43_P_NMU    32'h00000026
`define NOC2_XBR2X4__REG_HIGH_ID43_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID44_P_NMU    32'h00000027
`define NOC2_XBR2X4__REG_HIGH_ID44_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID45_P_NMU    32'h00000028
`define NOC2_XBR2X4__REG_HIGH_ID45_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID46_P_NMU    32'h00000029
`define NOC2_XBR2X4__REG_HIGH_ID46_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID47_P_NMU    32'h0000002a
`define NOC2_XBR2X4__REG_HIGH_ID47_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID48_P_NMU    32'h0000002b
`define NOC2_XBR2X4__REG_HIGH_ID48_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID49_P_NMU    32'h0000002c
`define NOC2_XBR2X4__REG_HIGH_ID49_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID4_P_NMU    32'h0000002d
`define NOC2_XBR2X4__REG_HIGH_ID4_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID50_P_NMU    32'h0000002e
`define NOC2_XBR2X4__REG_HIGH_ID50_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID51_P_NMU    32'h0000002f
`define NOC2_XBR2X4__REG_HIGH_ID51_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID52_P_NMU    32'h00000030
`define NOC2_XBR2X4__REG_HIGH_ID52_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID53_P_NMU    32'h00000031
`define NOC2_XBR2X4__REG_HIGH_ID53_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID54_P_NMU    32'h00000032
`define NOC2_XBR2X4__REG_HIGH_ID54_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID55_P_NMU    32'h00000033
`define NOC2_XBR2X4__REG_HIGH_ID55_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID56_P_NMU    32'h00000034
`define NOC2_XBR2X4__REG_HIGH_ID56_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID57_P_NMU    32'h00000035
`define NOC2_XBR2X4__REG_HIGH_ID57_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID58_P_NMU    32'h00000036
`define NOC2_XBR2X4__REG_HIGH_ID58_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID59_P_NMU    32'h00000037
`define NOC2_XBR2X4__REG_HIGH_ID59_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID5_P_NMU    32'h00000038
`define NOC2_XBR2X4__REG_HIGH_ID5_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID60_P_NMU    32'h00000039
`define NOC2_XBR2X4__REG_HIGH_ID60_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID61_P_NMU    32'h0000003a
`define NOC2_XBR2X4__REG_HIGH_ID61_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID62_P_NMU    32'h0000003b
`define NOC2_XBR2X4__REG_HIGH_ID62_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID63_P_NMU    32'h0000003c
`define NOC2_XBR2X4__REG_HIGH_ID63_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID6_P_NMU    32'h0000003d
`define NOC2_XBR2X4__REG_HIGH_ID6_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID7_P_NMU    32'h0000003e
`define NOC2_XBR2X4__REG_HIGH_ID7_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID8_P_NMU    32'h0000003f
`define NOC2_XBR2X4__REG_HIGH_ID8_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_HIGH_ID9_P_NMU    32'h00000040
`define NOC2_XBR2X4__REG_HIGH_ID9_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_ID    32'h00000041
`define NOC2_XBR2X4__REG_ID_SZ 10

`define NOC2_XBR2X4__REG_LOW_ID0_P_NMU    32'h00000042
`define NOC2_XBR2X4__REG_LOW_ID0_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID10_P_NMU    32'h00000043
`define NOC2_XBR2X4__REG_LOW_ID10_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID11_P_NMU    32'h00000044
`define NOC2_XBR2X4__REG_LOW_ID11_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID12_P_NMU    32'h00000045
`define NOC2_XBR2X4__REG_LOW_ID12_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID13_P_NMU    32'h00000046
`define NOC2_XBR2X4__REG_LOW_ID13_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID14_P_NMU    32'h00000047
`define NOC2_XBR2X4__REG_LOW_ID14_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID15_P_NMU    32'h00000048
`define NOC2_XBR2X4__REG_LOW_ID15_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID1_P_NMU    32'h00000049
`define NOC2_XBR2X4__REG_LOW_ID1_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID2_P_NMU    32'h0000004a
`define NOC2_XBR2X4__REG_LOW_ID2_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID3_P_NMU    32'h0000004b
`define NOC2_XBR2X4__REG_LOW_ID3_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID4_P_NMU    32'h0000004c
`define NOC2_XBR2X4__REG_LOW_ID4_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID5_P_NMU    32'h0000004d
`define NOC2_XBR2X4__REG_LOW_ID5_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID6_P_NMU    32'h0000004e
`define NOC2_XBR2X4__REG_LOW_ID6_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID7_P_NMU    32'h0000004f
`define NOC2_XBR2X4__REG_LOW_ID7_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID8_P_NMU    32'h00000050
`define NOC2_XBR2X4__REG_LOW_ID8_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_LOW_ID9_P_NMU    32'h00000051
`define NOC2_XBR2X4__REG_LOW_ID9_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_MID_ID0_P_NMU    32'h00000052
`define NOC2_XBR2X4__REG_MID_ID0_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_MID_ID1_P_NMU    32'h00000053
`define NOC2_XBR2X4__REG_MID_ID1_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_MID_ID2_P_NMU    32'h00000054
`define NOC2_XBR2X4__REG_MID_ID2_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_MID_ID3_P_NMU    32'h00000055
`define NOC2_XBR2X4__REG_MID_ID3_P_NMU_SZ 12

`define NOC2_XBR2X4__REG_NOC_CTL    32'h00000056
`define NOC2_XBR2X4__REG_NOC_CTL_SZ 16

`define NOC2_XBR2X4__REG_P00_P_NMU_0_VCA_TOKEN    32'h00000057
`define NOC2_XBR2X4__REG_P00_P_NMU_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P00_P_NMU_1_VCA_TOKEN    32'h00000058
`define NOC2_XBR2X4__REG_P00_P_NMU_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P01_P_NSU_0_VCA_TOKEN    32'h00000059
`define NOC2_XBR2X4__REG_P01_P_NSU_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P01_P_NSU_1_VCA_TOKEN    32'h0000005a
`define NOC2_XBR2X4__REG_P01_P_NSU_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P10_P_NMU_0_VCA_TOKEN    32'h0000005b
`define NOC2_XBR2X4__REG_P10_P_NMU_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P10_P_NMU_1_VCA_TOKEN    32'h0000005c
`define NOC2_XBR2X4__REG_P10_P_NMU_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P11_P_NSU_0_VCA_TOKEN    32'h0000005d
`define NOC2_XBR2X4__REG_P11_P_NSU_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P11_P_NSU_1_VCA_TOKEN    32'h0000005e
`define NOC2_XBR2X4__REG_P11_P_NSU_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P20_P_NMU_0_VCA_TOKEN    32'h0000005f
`define NOC2_XBR2X4__REG_P20_P_NMU_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P20_P_NMU_1_VCA_TOKEN    32'h00000060
`define NOC2_XBR2X4__REG_P20_P_NMU_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P21_P_NSU_0_VCA_TOKEN    32'h00000061
`define NOC2_XBR2X4__REG_P21_P_NSU_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P21_P_NSU_1_VCA_TOKEN    32'h00000062
`define NOC2_XBR2X4__REG_P21_P_NSU_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P30_P_NMU_0_VCA_TOKEN    32'h00000063
`define NOC2_XBR2X4__REG_P30_P_NMU_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P30_P_NMU_1_VCA_TOKEN    32'h00000064
`define NOC2_XBR2X4__REG_P30_P_NMU_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P31_P_NSU_0_VCA_TOKEN    32'h00000065
`define NOC2_XBR2X4__REG_P31_P_NSU_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P31_P_NSU_1_VCA_TOKEN    32'h00000066
`define NOC2_XBR2X4__REG_P31_P_NSU_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU0_P0_0_VCA_TOKEN    32'h00000067
`define NOC2_XBR2X4__REG_P_NMU0_P0_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU0_P0_1_VCA_TOKEN    32'h00000068
`define NOC2_XBR2X4__REG_P_NMU0_P0_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU1_P1_0_VCA_TOKEN    32'h00000069
`define NOC2_XBR2X4__REG_P_NMU1_P1_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU1_P1_1_VCA_TOKEN    32'h0000006a
`define NOC2_XBR2X4__REG_P_NMU1_P1_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU2_P2_0_VCA_TOKEN    32'h0000006b
`define NOC2_XBR2X4__REG_P_NMU2_P2_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU2_P2_1_VCA_TOKEN    32'h0000006c
`define NOC2_XBR2X4__REG_P_NMU2_P2_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU3_P3_0_VCA_TOKEN    32'h0000006d
`define NOC2_XBR2X4__REG_P_NMU3_P3_0_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NMU3_P3_1_VCA_TOKEN    32'h0000006e
`define NOC2_XBR2X4__REG_P_NMU3_P3_1_VCA_TOKEN_SZ 32

`define NOC2_XBR2X4__REG_P_NSU0_P0_0_VCA_TOKEN    32'h0000006f
`define NOC2_XBR2X4__REG_P_NSU0_P0_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU0_P0_1_VCA_TOKEN    32'h00000070
`define NOC2_XBR2X4__REG_P_NSU0_P0_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU1_P1_0_VCA_TOKEN    32'h00000071
`define NOC2_XBR2X4__REG_P_NSU1_P1_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU1_P1_1_VCA_TOKEN    32'h00000072
`define NOC2_XBR2X4__REG_P_NSU1_P1_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU2_P2_0_VCA_TOKEN    32'h00000073
`define NOC2_XBR2X4__REG_P_NSU2_P2_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU2_P2_1_VCA_TOKEN    32'h00000074
`define NOC2_XBR2X4__REG_P_NSU2_P2_1_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU3_P3_0_VCA_TOKEN    32'h00000075
`define NOC2_XBR2X4__REG_P_NSU3_P3_0_VCA_TOKEN_SZ 16

`define NOC2_XBR2X4__REG_P_NSU3_P3_1_VCA_TOKEN    32'h00000076
`define NOC2_XBR2X4__REG_P_NSU3_P3_1_VCA_TOKEN_SZ 16

`endif  // B_NOC2_XBR2X4_DEFINES_VH