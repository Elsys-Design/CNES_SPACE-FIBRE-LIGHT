`include "B_IBUFDS_INTERMDISABLE_defines.vh"

reg [`IBUFDS_INTERMDISABLE_DATA_SZ-1:0] ATTR [0:`IBUFDS_INTERMDISABLE_ADDR_N-1];
reg [`IBUFDS_INTERMDISABLE__DIFF_TERM_SZ:1] DIFF_TERM_REG = DIFF_TERM;
reg [`IBUFDS_INTERMDISABLE__DQS_BIAS_SZ:1] DQS_BIAS_REG = DQS_BIAS;
reg [`IBUFDS_INTERMDISABLE__IBUF_LOW_PWR_SZ:1] IBUF_LOW_PWR_REG = IBUF_LOW_PWR;
reg [`IBUFDS_INTERMDISABLE__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IBUFDS_INTERMDISABLE__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`IBUFDS_INTERMDISABLE__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IBUFDS_INTERMDISABLE__DIFF_TERM] = DIFF_TERM;
  ATTR[`IBUFDS_INTERMDISABLE__DQS_BIAS] = DQS_BIAS;
  ATTR[`IBUFDS_INTERMDISABLE__IBUF_LOW_PWR] = IBUF_LOW_PWR;
  ATTR[`IBUFDS_INTERMDISABLE__IOSTANDARD] = IOSTANDARD;
  ATTR[`IBUFDS_INTERMDISABLE__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`IBUFDS_INTERMDISABLE__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  DIFF_TERM_REG = ATTR[`IBUFDS_INTERMDISABLE__DIFF_TERM];
  DQS_BIAS_REG = ATTR[`IBUFDS_INTERMDISABLE__DQS_BIAS];
  IBUF_LOW_PWR_REG = ATTR[`IBUFDS_INTERMDISABLE__IBUF_LOW_PWR];
  IOSTANDARD_REG = ATTR[`IBUFDS_INTERMDISABLE__IOSTANDARD];
  SIM_DEVICE_REG = ATTR[`IBUFDS_INTERMDISABLE__SIM_DEVICE];
  USE_IBUFDISABLE_REG = ATTR[`IBUFDS_INTERMDISABLE__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IBUFDS_INTERMDISABLE_ADDR_SZ-1:0] addr;
  input  [`IBUFDS_INTERMDISABLE_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IBUFDS_INTERMDISABLE_DATA_SZ-1:0] read_attr;
  input  [`IBUFDS_INTERMDISABLE_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
