// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HPLL_DEFINES_VH
`else
`define B_HPLL_DEFINES_VH

// Look-up table parameters
//

`define HPLL_ADDR_N  49
`define HPLL_ADDR_SZ 32
`define HPLL_DATA_SZ 64

// Attribute addresses
//

`define HPLL__CLKFBOUT_MULT    32'h00000000
`define HPLL__CLKFBOUT_MULT_SZ 32

`define HPLL__CLKFBOUT_PHASE    32'h00000001
`define HPLL__CLKFBOUT_PHASE_SZ 64

`define HPLL__CLKIN_FREQ_MAX    32'h00000002
`define HPLL__CLKIN_FREQ_MAX_SZ 64

`define HPLL__CLKIN_FREQ_MIN    32'h00000003
`define HPLL__CLKIN_FREQ_MIN_SZ 64

`define HPLL__CLKIN_PERIOD    32'h00000004
`define HPLL__CLKIN_PERIOD_SZ 64

`define HPLL__CLKOUT0_DIVIDE    32'h00000005
`define HPLL__CLKOUT0_DIVIDE_SZ 32

`define HPLL__CLKOUT0_DUTY_CYCLE    32'h00000006
`define HPLL__CLKOUT0_DUTY_CYCLE_SZ 64

`define HPLL__CLKOUT0_PHASE    32'h00000007
`define HPLL__CLKOUT0_PHASE_SZ 64

`define HPLL__CLKOUT0_PHASE_CTRL    32'h00000008
`define HPLL__CLKOUT0_PHASE_CTRL_SZ 2

`define HPLL__CLKOUT1_DIVIDE    32'h00000009
`define HPLL__CLKOUT1_DIVIDE_SZ 32

`define HPLL__CLKOUT1_DUTY_CYCLE    32'h0000000a
`define HPLL__CLKOUT1_DUTY_CYCLE_SZ 64

`define HPLL__CLKOUT1_PHASE    32'h0000000b
`define HPLL__CLKOUT1_PHASE_SZ 64

`define HPLL__CLKOUT1_PHASE_CTRL    32'h0000000c
`define HPLL__CLKOUT1_PHASE_CTRL_SZ 2

`define HPLL__CLKOUT2_DIVIDE    32'h0000000d
`define HPLL__CLKOUT2_DIVIDE_SZ 32

`define HPLL__CLKOUT2_DUTY_CYCLE    32'h0000000e
`define HPLL__CLKOUT2_DUTY_CYCLE_SZ 64

`define HPLL__CLKOUT2_PHASE    32'h0000000f
`define HPLL__CLKOUT2_PHASE_SZ 64

`define HPLL__CLKOUT2_PHASE_CTRL    32'h00000010
`define HPLL__CLKOUT2_PHASE_CTRL_SZ 2

`define HPLL__CLKOUT3_DIVIDE    32'h00000011
`define HPLL__CLKOUT3_DIVIDE_SZ 32

`define HPLL__CLKOUT3_DUTY_CYCLE    32'h00000012
`define HPLL__CLKOUT3_DUTY_CYCLE_SZ 64

`define HPLL__CLKOUT3_PHASE    32'h00000013
`define HPLL__CLKOUT3_PHASE_SZ 64

`define HPLL__CLKOUT3_PHASE_CTRL    32'h00000014
`define HPLL__CLKOUT3_PHASE_CTRL_SZ 2

`define HPLL__CLKOUTPHY_CASCIN_EN    32'h00000015
`define HPLL__CLKOUTPHY_CASCIN_EN_SZ 1

`define HPLL__CLKOUTPHY_CASCOUT_EN    32'h00000016
`define HPLL__CLKOUTPHY_CASCOUT_EN_SZ 1

`define HPLL__CLKOUTPHY_DIVIDE    32'h00000017
`define HPLL__CLKOUTPHY_DIVIDE_SZ 40

`define HPLL__CLKPFD_FREQ_MAX    32'h00000018
`define HPLL__CLKPFD_FREQ_MAX_SZ 64

`define HPLL__CLKPFD_FREQ_MIN    32'h00000019
`define HPLL__CLKPFD_FREQ_MIN_SZ 64

`define HPLL__DESKEW2_MUXIN_SEL    32'h0000001a
`define HPLL__DESKEW2_MUXIN_SEL_SZ 1

`define HPLL__DESKEW_DELAY1    32'h0000001b
`define HPLL__DESKEW_DELAY1_SZ 32

`define HPLL__DESKEW_DELAY2    32'h0000001c
`define HPLL__DESKEW_DELAY2_SZ 32

`define HPLL__DESKEW_DELAY_EN1    32'h0000001d
`define HPLL__DESKEW_DELAY_EN1_SZ 40

`define HPLL__DESKEW_DELAY_EN2    32'h0000001e
`define HPLL__DESKEW_DELAY_EN2_SZ 40

`define HPLL__DESKEW_DELAY_PATH1    32'h0000001f
`define HPLL__DESKEW_DELAY_PATH1_SZ 40

`define HPLL__DESKEW_DELAY_PATH2    32'h00000020
`define HPLL__DESKEW_DELAY_PATH2_SZ 40

`define HPLL__DESKEW_MUXIN_SEL    32'h00000021
`define HPLL__DESKEW_MUXIN_SEL_SZ 1

`define HPLL__DIV4_CLKOUT012    32'h00000022
`define HPLL__DIV4_CLKOUT012_SZ 1

`define HPLL__DIV4_CLKOUT3    32'h00000023
`define HPLL__DIV4_CLKOUT3_SZ 1

`define HPLL__DIVCLK_DIVIDE    32'h00000024
`define HPLL__DIVCLK_DIVIDE_SZ 32

`define HPLL__IS_CLKFB1_DESKEW_INVERTED    32'h00000025
`define HPLL__IS_CLKFB1_DESKEW_INVERTED_SZ 1

`define HPLL__IS_CLKFB2_DESKEW_INVERTED    32'h00000026
`define HPLL__IS_CLKFB2_DESKEW_INVERTED_SZ 1

`define HPLL__IS_CLKIN1_DESKEW_INVERTED    32'h00000027
`define HPLL__IS_CLKIN1_DESKEW_INVERTED_SZ 1

`define HPLL__IS_CLKIN2_DESKEW_INVERTED    32'h00000028
`define HPLL__IS_CLKIN2_DESKEW_INVERTED_SZ 1

`define HPLL__IS_CLKIN_INVERTED    32'h00000029
`define HPLL__IS_CLKIN_INVERTED_SZ 1

`define HPLL__IS_PSEN_INVERTED    32'h0000002a
`define HPLL__IS_PSEN_INVERTED_SZ 1

`define HPLL__IS_PSINCDEC_INVERTED    32'h0000002b
`define HPLL__IS_PSINCDEC_INVERTED_SZ 1

`define HPLL__IS_PWRDWN_INVERTED    32'h0000002c
`define HPLL__IS_PWRDWN_INVERTED_SZ 1

`define HPLL__IS_RST_INVERTED    32'h0000002d
`define HPLL__IS_RST_INVERTED_SZ 1

`define HPLL__REF_JITTER    32'h0000002e
`define HPLL__REF_JITTER_SZ 64

`define HPLL__VCOCLK_FREQ_MAX    32'h0000002f
`define HPLL__VCOCLK_FREQ_MAX_SZ 64

`define HPLL__VCOCLK_FREQ_MIN    32'h00000030
`define HPLL__VCOCLK_FREQ_MIN_SZ 64

`endif  // B_HPLL_DEFINES_VH