// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC2_NSU128_DEFINES_VH
`else
`define B_NOC2_NSU128_DEFINES_VH

// Look-up table parameters
//

`define NOC2_NSU128_ADDR_N  40
`define NOC2_NSU128_ADDR_SZ 32
`define NOC2_NSU128_DATA_SZ 12

// Attribute addresses
//

`define NOC2_NSU128__REG_AFWM_EN    32'h00000000
`define NOC2_NSU128__REG_AFWM_EN_SZ 1

`define NOC2_NSU128__REG_AFWM_INTR_EN    32'h00000001
`define NOC2_NSU128__REG_AFWM_INTR_EN_SZ 1

`define NOC2_NSU128__REG_AFWM_TIMEOUT_ERR_EN    32'h00000002
`define NOC2_NSU128__REG_AFWM_TIMEOUT_ERR_EN_SZ 5

`define NOC2_NSU128__REG_AXI_LOOPBACK    32'h00000003
`define NOC2_NSU128__REG_AXI_LOOPBACK_SZ 2

`define NOC2_NSU128__REG_COMP_ID_INDEX0    32'h00000004
`define NOC2_NSU128__REG_COMP_ID_INDEX0_SZ 5

`define NOC2_NSU128__REG_COMP_ID_INDEX1    32'h00000005
`define NOC2_NSU128__REG_COMP_ID_INDEX1_SZ 5

`define NOC2_NSU128__REG_COMP_ID_MODE    32'h00000006
`define NOC2_NSU128__REG_COMP_ID_MODE_SZ 1

`define NOC2_NSU128__REG_DISABLE_EX_MON    32'h00000007
`define NOC2_NSU128__REG_DISABLE_EX_MON_SZ 1

`define NOC2_NSU128__REG_DST_ID_MASK    32'h00000008
`define NOC2_NSU128__REG_DST_ID_MASK_SZ 12

`define NOC2_NSU128__REG_DWIDTH    32'h00000009
`define NOC2_NSU128__REG_DWIDTH_SZ 3

`define NOC2_NSU128__REG_ECC_CHK_EN    32'h0000000a
`define NOC2_NSU128__REG_ECC_CHK_EN_SZ 1

`define NOC2_NSU128__REG_FIXED_COMP_ID    32'h0000000b
`define NOC2_NSU128__REG_FIXED_COMP_ID_SZ 2

`define NOC2_NSU128__REG_MODE_SELECT    32'h0000000c
`define NOC2_NSU128__REG_MODE_SELECT_SZ 2

`define NOC2_NSU128__REG_ODISABLE_AXI_RESP    32'h0000000d
`define NOC2_NSU128__REG_ODISABLE_AXI_RESP_SZ 1

`define NOC2_NSU128__REG_OUTSTANDING_RD_TXN    32'h0000000e
`define NOC2_NSU128__REG_OUTSTANDING_RD_TXN_SZ 6

`define NOC2_NSU128__REG_OUTSTANDING_WR_TXN    32'h0000000f
`define NOC2_NSU128__REG_OUTSTANDING_WR_TXN_SZ 6

`define NOC2_NSU128__REG_PAR_CHK    32'h00000010
`define NOC2_NSU128__REG_PAR_CHK_SZ 2

`define NOC2_NSU128__REG_RDTRK_VCA_TOKEN0    32'h00000011
`define NOC2_NSU128__REG_RDTRK_VCA_TOKEN0_SZ 8

`define NOC2_NSU128__REG_RDTRK_VCA_TOKEN1    32'h00000012
`define NOC2_NSU128__REG_RDTRK_VCA_TOKEN1_SZ 8

`define NOC2_NSU128__REG_RD_REQ_VC_MAP0    32'h00000013
`define NOC2_NSU128__REG_RD_REQ_VC_MAP0_SZ 3

`define NOC2_NSU128__REG_RD_REQ_VC_MAP1    32'h00000014
`define NOC2_NSU128__REG_RD_REQ_VC_MAP1_SZ 3

`define NOC2_NSU128__REG_RD_RESP_VC_MAP0    32'h00000015
`define NOC2_NSU128__REG_RD_RESP_VC_MAP0_SZ 3

`define NOC2_NSU128__REG_RD_RESP_VC_MAP1    32'h00000016
`define NOC2_NSU128__REG_RD_RESP_VC_MAP1_SZ 3

`define NOC2_NSU128__REG_RD_VCA_TOKEN0    32'h00000017
`define NOC2_NSU128__REG_RD_VCA_TOKEN0_SZ 8

`define NOC2_NSU128__REG_RD_VCA_TOKEN1    32'h00000018
`define NOC2_NSU128__REG_RD_VCA_TOKEN1_SZ 8

`define NOC2_NSU128__REG_SRC    32'h00000019
`define NOC2_NSU128__REG_SRC_SZ 12

`define NOC2_NSU128__REG_TBASE_AXI_TIMEOUT    32'h0000001a
`define NOC2_NSU128__REG_TBASE_AXI_TIMEOUT_SZ 4

`define NOC2_NSU128__REG_TBASE_TRK_TIMEOUT    32'h0000001b
`define NOC2_NSU128__REG_TBASE_TRK_TIMEOUT_SZ 4

`define NOC2_NSU128__REG_VMAP_OUT_RD_TOKEN0    32'h0000001c
`define NOC2_NSU128__REG_VMAP_OUT_RD_TOKEN0_SZ 8

`define NOC2_NSU128__REG_VMAP_OUT_RD_TOKEN1    32'h0000001d
`define NOC2_NSU128__REG_VMAP_OUT_RD_TOKEN1_SZ 8

`define NOC2_NSU128__REG_VMAP_OUT_WR_TOKEN0    32'h0000001e
`define NOC2_NSU128__REG_VMAP_OUT_WR_TOKEN0_SZ 8

`define NOC2_NSU128__REG_VMAP_OUT_WR_TOKEN1    32'h0000001f
`define NOC2_NSU128__REG_VMAP_OUT_WR_TOKEN1_SZ 8

`define NOC2_NSU128__REG_WRTRK_VCA_TOKEN0    32'h00000020
`define NOC2_NSU128__REG_WRTRK_VCA_TOKEN0_SZ 8

`define NOC2_NSU128__REG_WRTRK_VCA_TOKEN1    32'h00000021
`define NOC2_NSU128__REG_WRTRK_VCA_TOKEN1_SZ 8

`define NOC2_NSU128__REG_WR_REQ_VC_MAP0    32'h00000022
`define NOC2_NSU128__REG_WR_REQ_VC_MAP0_SZ 3

`define NOC2_NSU128__REG_WR_REQ_VC_MAP1    32'h00000023
`define NOC2_NSU128__REG_WR_REQ_VC_MAP1_SZ 3

`define NOC2_NSU128__REG_WR_RESP_VC_MAP0    32'h00000024
`define NOC2_NSU128__REG_WR_RESP_VC_MAP0_SZ 3

`define NOC2_NSU128__REG_WR_RESP_VC_MAP1    32'h00000025
`define NOC2_NSU128__REG_WR_RESP_VC_MAP1_SZ 3

`define NOC2_NSU128__REG_WR_VCA_TOKEN0    32'h00000026
`define NOC2_NSU128__REG_WR_VCA_TOKEN0_SZ 8

`define NOC2_NSU128__REG_WR_VCA_TOKEN1    32'h00000027
`define NOC2_NSU128__REG_WR_VCA_TOKEN1_SZ 8

`endif  // B_NOC2_NSU128_DEFINES_VH