library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.data_link_lib.all;

entity subpart_tb is
end subpart_tb;

architecture Behavioral of subpart_tb is
  -- Déclaration des composants
  COMPONENT data_encpasulation IS
    GENERIC (
        G_VC_NUM                       : INTEGER := 8                                                  --! Number of virtual channel
    );
    PORT (
      RST_N                            : IN  std_logic;                                    --! global reset
      CLK                              : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DMAC interface
      DATA_DMAC                        : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      NEW_WORD_DMAC                    : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      NEW_PACKET_DMAC                  : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      END_PACKET_DMAC                  : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      TYPE_FRAME_DMAC                  : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);                 --! Flag EMPTY of the FIFO RX
      VIRTUAL_CHANNEL_DMAC             : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_TYPE_DMAC                     : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_CHANNEL_DMAC                  : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      BC_STATUS_DMAC                    : in std_logic_vector (2-1 downto 0);
      MULT_CHANNEL_DMAC                : IN std_logic_vector (G_VC_NUM-1 DOWNTO 0);
      -- DSCOM interface
      NEW_WORD_DENC                    : OUT  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DENC                        : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DENC              : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DENC                  : OUT  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);                 --! Flag EMPTY of the FIFO RX
      END_FRAME_DENC                   : OUT  std_logic
    );
  END COMPONENT;

  COMPONENT data_seq_compute IS
    PORT (
      RST_N                 : IN  std_logic;                                    --! global reset
      CLK                   : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DENC interface
      NEW_WORD_DENC         : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DENC        : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DENC   : IN  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DENC       : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DENC        : IN  std_logic;
      -- DCCOM interface
      NEW_WORD_DSCOM        : OUT  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DSCOM       : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DSCOM  : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DSCOM      : OUT  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DSCOM       : OUT  std_logic
    );
  END COMPONENT;

  COMPONENT data_crc_compute IS
    PORT (
      RST_N                 : IN  std_logic;                                    --! global reset
      CLK                   : IN  std_logic;                                    --! Clock generated by GTY IP
      -- DSCOM interface
      NEW_WORD_DSCOM        : IN  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
      DATA_DSCOM            : IN  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);   --! Data parallel from Lane Layer
      VALID_K_CHARAC_DSCOM  : IN  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      TYPE_FRAME_DSCOM      : IN  std_logic_vector(C_TYPE_FRAME_LENGTH-1 DOWNTO 0);
      END_FRAME_DSCOM       : IN  std_logic;
      -- FIFO_TX_LANE interface
      FIFO_FULL_TX_LANE     : IN  std_logic;
      VALID_K_CHARAC_DCCOM  : OUT  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 DOWNTO 0);
      DATA_DCCOM            : OUT  std_logic_vector(C_DATA_LENGTH-1 DOWNTO 0);    -- Data write bus
      NEW_WORD_DCCOM        : OUT  std_logic                                -- Write command
    );
  END COMPONENT;

  COMPONENT data_word_id_fsm IS
  port (
    RST_N                   : in  std_logic;                                    --! global reset
    CLK                     : in  std_logic;                                    --! Clock generated by GTY IP
    LINK_RESET              : in  std_logic;                                    --! Link Reset command 
    -- PHY PLUS LANE layer interface
    FIFO_RX_DATA_VALID_PPL  : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    FIFO_RX_RD_EN_PPL       : out  std_logic;                                   --! Flag to read data in FIFO RX  
    DATA_RX_PPL             : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    VALID_K_CHARAC_PPL    : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);               --! K charachter valid in the 32-bit DATA_RX_PPL vector
    -- DCCHECK layer interface
    TYPE_FRAME_DWI          : out  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    NEW_WORD_DWI            : out   std_logic;   
    END_FRAME_DWI           : out  std_logic;
    DATA_DWI                : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    SEQ_NUM_DWI             : out  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX 
    CRC_16B_DWI             : out  std_logic_vector(15 downto 0);                --! Flag EMPTY of the FIFO RX
    CRC_8B_DWI              : out  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
    -- OTHER
    CRC_ERR                 : in   std_logic;   
    SEQ_ERR                 : in   std_logic;   
    FRAME_ERR               : out   std_logic  
  );
  END COMPONENT;

  COMPONENT data_CRC_check IS
  port(
    RST_N              : in  std_logic;                                    --! global reset
    CLK                : in  std_logic;                                    --! Clock generated by GTY IP
    -- DWI interface
    DATA_DWI           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    NEW_WORD_DWI       : in  std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    END_FRAME_DWI      : in  std_logic;
    SEQ_NUM_DWI        : in  std_logic_vector(7 downto 0);
    CRC_16B_DWI        : in  std_logic_vector(15 downto 0);                --! Flag EMPTY of the FIFO RX
    CRC_8B_DWI         : in  std_logic_vector(7 downto 0);                 --! Flag EMPTY of the FIFO RX
    TYPE_FRAME_DWI     : in  std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);                 --! Flag EMPTY of the FIFO RX
    -- DWI interface
    NEW_WORD_DCCHECK   : out std_logic;                                    --! Flag DATA_VALID of the FIFO RX from Lane layer
    DATA_DCCHECK       : out std_logic_vector(C_DATA_LENGTH-1 downto 0);   --! Data parallel from Lane Layer
    END_FRAME_DCCHECK  : out std_logic;
    TYPE_FRAME_DCCHECK : out std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);                 --! Flag EMPTY of the FIFO RX
    SEQ_NUM_DCCHECK    : out std_logic_vector(7 downto 0);
    CRC_ERR            : out std_logic

  );
  END COMPONENT;

  COMPONENT data_seq_check IS
  port (
    RST_N                  : in  std_logic;                                    --! global reset
    CLK                    : in  std_logic;                                    --! Clock generated by GTY IP
    -- DCCHECK interface
    DATA_DCCHECK           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);                   --! Data parallel from Lane Layer
    SEQ_NUM_DCCHECK        : in  STD_LOGIC_VECTOR(7 downto 0);                      --! Flag EMPTY of the FIFO RX
    END_FRAME_DCCHECK      : in std_logic;
    REC_POLARITY_FLG       : in  std_logic;                                         --! Flag EMPTY of the FIFO RX
    TYPE_FRAME_DCCHECK     : in  STD_LOGIC_VECTOR(C_TYPE_FRAME_LENGTH-1 downto 0);  --! Flag EMPTY of the FIFO RX
    NEW_WORD_DCCHECK       : in  std_logic;  
    -- FIFO signals
    DATA_DSCHECK           : out  std_logic_vector(C_DATA_LENGTH-1 downto 0);    -- Data write bus
    NEW_WORD_DSCHECK       : out  std_logic;                                -- Write command
    END_FRAME_DSCHECK      : out std_logic;
    SEQ_NUM_ERR            : out std_logic;
    FIFO_FULL              : in std_logic 
  );
  END COMPONENT;

    -- Constants
    constant G_VC_NUM               : integer := 8;

    -- Clock and Reset
    signal CLK     : std_logic := '0';
    signal RST_N   : std_logic := '0';

    -- DMAC interface signals
    signal DATA_DMAC                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal NEW_WORD_DMAC             : std_logic;
    signal NEW_PACKET_DMAC           : std_logic;
    signal END_PACKET_DMAC           : std_logic;
    signal TYPE_FRAME_DMAC           : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    signal VIRTUAL_CHANNEL_DMAC      : std_logic_vector(G_VC_NUM-1 downto 0);
    signal BC_TYPE_DMAC              : std_logic_vector(G_VC_NUM-1 downto 0);
    signal BC_CHANNEL_DMAC           : std_logic_vector(G_VC_NUM-1 downto 0);
    signal BC_STATUS_DMAC            : std_logic_vector(2-1 downto 0);
    signal MULT_CHANNEL_DMAC         : std_logic_vector(G_VC_NUM-1 downto 0);

    -- DENC interface signals
    signal NEW_WORD_DENC             : std_logic;
    signal DATA_DENC                 : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal VALID_K_CHARAC_DENC       : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
    signal TYPE_FRAME_DENC           : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    signal END_FRAME_DENC            : std_logic;

    -- DSCOM interface signals
    signal NEW_WORD_DSCOM            : std_logic;
    signal DATA_DSCOM           : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal VALID_K_CHARAC_DSCOM      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
    signal TYPE_FRAME_DSCOM          : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    signal END_FRAME_DSCOM           : std_logic;

    -- FIFO_TX_LANE interface signals
    signal FIFO_FULL_TX_LANE         : std_logic:='0';
    signal VALID_K_CHARAC_DCCOM      : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
    signal DATA_DCCOM                : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal NEW_WORD_DCCOM            : std_logic;

    -- DWI interface signals
    signal DATA_DWI                  : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal NEW_WORD_DWI              : std_logic;
    signal END_FRAME_DWI              : std_logic;
    signal SEQ_NUM_DWI                : std_logic_vector(7 downto 0);
    signal CRC_16B_DWI               : std_logic_vector(15 downto 0);
    signal CRC_8B_DWI                : std_logic_vector(7 downto 0);
    signal TYPE_FRAME_DWI            : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);

    -- CRC Check signals
    signal NEW_WORD_DCCHECK          : std_logic;
    signal DATA_DCCHECK         : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal SEQ_NUM_DCCHECK           : std_logic_vector(7 downto 0);
    signal END_FRAME_DCCHECK            : std_logic;
    signal CRC_ERR                   : std_logic;

    -- Sequence Check signals
    signal REC_POLARITY_FLG          : std_logic;
    signal TYPE_FRAME_DCCHECK        : std_logic_vector(C_TYPE_FRAME_LENGTH-1 downto 0);
    signal SEQ_NUM_ERR               : std_logic;
    signal DATA_DSCHECK         : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal END_FRAME_DSCHECK               : std_logic;
    signal NEW_WORD_DSCHECK          : std_logic;
    signal FIFO_FULL                 : std_logic:='0';

    -- PHY PLUS LANE layer interface signals
    signal FIFO_RX_DATA_VALID_PPL    : std_logic;
    signal FIFO_RX_RD_EN_PPL         : std_logic;
    signal DATA_RX_PPL               : std_logic_vector(C_DATA_LENGTH-1 downto 0);
    signal VALID_K_CHARAC_RX_PPL     : std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);
    signal LINK_RESET                : std_logic;
    signal FRAME_ERR                 : std_logic;
    signal SEQ_ERR                    : std_logic;

    -- Clock process definitions
    constant CLOCK_PERIOD : time := 10 ns;
begin

    -- Clock process
    CLK_process :process
    begin
        CLK <= '0';
        wait for CLOCK_PERIOD/2;
        CLK <= '1';
        wait for CLOCK_PERIOD/2;
    end process;

    main_process: process
    begin
      RST_N <= '0';
      wait for 20 ns;
      RST_N          <= '1';
      wait for CLOCK_PERIOD/2;
      DATA_DMAC            <=(others =>'0');  
      NEW_WORD_DMAC        <= '0';
      NEW_PACKET_DMAC      <= '0';
      END_PACKET_DMAC      <= '0';
      TYPE_FRAME_DMAC      <=(others =>'0');  
      VIRTUAL_CHANNEL_DMAC <=(others =>'0');  
      BC_TYPE_DMAC         <=(others =>'0');  
      BC_CHANNEL_DMAC      <=(others =>'0');    
      MULT_CHANNEL_DMAC    <=(others =>'0');   

      wait for 2 * CLOCK_PERIOD;
      TYPE_FRAME_DMAC      <= C_DATA_FRM;
      VIRTUAL_CHANNEL_DMAC <= std_logic_vector(to_unsigned(2,VIRTUAL_CHANNEL_DMAC'length));
      NEW_PACKET_DMAC      <= '1';

      wait for CLOCK_PERIOD;

      NEW_PACKET_DMAC      <= '0';
      END_PACKET_DMAC      <= '0';
      NEW_WORD_DMAC        <= '1';
      DATA_DMAC            <= C_RESERVED_SYMB & C_RESERVED_SYMB & C_RESERVED_SYMB & C_RESERVED_SYMB;

      wait for CLOCK_PERIOD;

      NEW_PACKET_DMAC      <= '0';
      END_PACKET_DMAC      <= '1';
      NEW_WORD_DMAC        <= '1';
      DATA_DMAC            <= C_FILL_SYMB & C_FILL_SYMB & C_FILL_SYMB& C_EOP_SYMB;

      wait for CLOCK_PERIOD;
      NEW_PACKET_DMAC      <= '0';
      END_PACKET_DMAC      <= '0';
      NEW_WORD_DMAC        <= '0';
      wait for CLOCK_PERIOD;
      DATA_DMAC            <= (others =>'0');  
      NEW_WORD_DMAC        <= '0';
      NEW_PACKET_DMAC      <= '0';
      END_PACKET_DMAC      <= '0';
      TYPE_FRAME_DMAC      <= (others =>'0');  
      VIRTUAL_CHANNEL_DMAC <= (others =>'0');  
      BC_TYPE_DMAC         <= (others =>'0');  
      BC_CHANNEL_DMAC      <= (others =>'0');    
      MULT_CHANNEL_DMAC    <= (others =>'0');   
      wait for CLOCK_PERIOD;
      wait;
    end process;

    -- Instantiate components
    UUT_data_encpasulation: entity work.data_encpasulation
        generic map (
            G_VC_NUM => G_VC_NUM
        )
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            DATA_DMAC             => DATA_DMAC,
            NEW_WORD_DMAC         => NEW_WORD_DMAC,
            NEW_PACKET_DMAC       => NEW_PACKET_DMAC,
            END_PACKET_DMAC       => END_PACKET_DMAC,
            TYPE_FRAME_DMAC       => TYPE_FRAME_DMAC,
            VIRTUAL_CHANNEL_DMAC  => VIRTUAL_CHANNEL_DMAC,
            BC_TYPE_DMAC          => BC_TYPE_DMAC,
            BC_CHANNEL_DMAC       => BC_CHANNEL_DMAC,
            BC_STATUS_DMAC        => BC_STATUS_DMAC,
            MULT_CHANNEL_DMAC     => MULT_CHANNEL_DMAC,
            NEW_WORD_DENC         => NEW_WORD_DENC,
            DATA_DENC             => DATA_DENC,
            VALID_K_CHARAC_DENC   => VALID_K_CHARAC_DENC,
            TYPE_FRAME_DENC       => TYPE_FRAME_DENC,
            END_FRAME_DENC        => END_FRAME_DENC
        );

    UUT_data_seq_compute: entity work.data_seq_compute
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            NEW_WORD_DENC         => NEW_WORD_DENC,
            DATA_DENC        => DATA_DENC,
            VALID_K_CHARAC_DENC   => VALID_K_CHARAC_DENC,
            TYPE_FRAME_DENC       => TYPE_FRAME_DENC,
            END_FRAME_DENC        => END_FRAME_DENC,
            NEW_WORD_DSCOM        => NEW_WORD_DSCOM,
            DATA_DSCOM       => DATA_DSCOM,
            VALID_K_CHARAC_DSCOM  => VALID_K_CHARAC_DSCOM,
            TYPE_FRAME_DSCOM      => TYPE_FRAME_DSCOM,
            END_FRAME_DSCOM       => END_FRAME_DSCOM
        );

    UUT_data_crc_compute: entity work.data_crc_compute
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            NEW_WORD_DSCOM        => NEW_WORD_DSCOM,
            DATA_DSCOM            => DATA_DSCOM,
            VALID_K_CHARAC_DSCOM  => VALID_K_CHARAC_DSCOM,
            TYPE_FRAME_DSCOM      => TYPE_FRAME_DSCOM,
            END_FRAME_DSCOM       => END_FRAME_DSCOM,
            FIFO_FULL_TX_LANE     => FIFO_FULL_TX_LANE,
            VALID_K_CHARAC_DCCOM  => VALID_K_CHARAC_DCCOM,
            DATA_DCCOM            => DATA_DCCOM,
            NEW_WORD_DCCOM        => NEW_WORD_DCCOM
        );

    UUT_data_word_id_fsm: entity work.data_word_id_fsm
        port map (
            RST_N                 => RST_N,
            CLK                   => CLK,
            LINK_RESET            => LINK_RESET,
            FIFO_RX_DATA_VALID_PPL=> NEW_WORD_DCCOM,
            FIFO_RX_RD_EN_PPL     => FIFO_RX_RD_EN_PPL,
            DATA_RX_PPL           => DATA_DCCOM,
            VALID_K_CHARAC_PPL  => VALID_K_CHARAC_DCCOM,
            TYPE_FRAME_DWI        => TYPE_FRAME_DWI,
            NEW_WORD_DWI          => NEW_WORD_DWI,
            END_FRAME_DWI         => END_FRAME_DWI,
            DATA_DWI              => DATA_DWI,
            SEQ_NUM_DWI           => SEQ_NUM_DWI,
            CRC_16B_DWI           => CRC_16B_DWI,
            CRC_8B_DWI            => CRC_8B_DWI,
            CRC_ERR               => CRC_ERR,
            SEQ_ERR               => SEQ_ERR,
            FRAME_ERR             => FRAME_ERR
        );

    UUT_data_CRC_check: entity work.data_CRC_check
        port map (
            RST_N              => RST_N,
            CLK                => CLK,
            DATA_DWI           => DATA_DWI,
            NEW_WORD_DWI       => NEW_WORD_DWI,
            END_FRAME_DWI         => END_FRAME_DWI,
            SEQ_NUM_DWI        => SEQ_NUM_DWI,
            CRC_16B_DWI        => CRC_16B_DWI,
            CRC_8B_DWI         => CRC_8B_DWI,
            TYPE_FRAME_DWI     => TYPE_FRAME_DWI,
            NEW_WORD_DCCHECK   => NEW_WORD_DCCHECK,
            DATA_DCCHECK  => DATA_DCCHECK,
            END_FRAME_DCCHECK         => END_FRAME_DCCHECK,
            TYPE_FRAME_DCCHECK     => TYPE_FRAME_DCCHECK,
            SEQ_NUM_DCCHECK    => SEQ_NUM_DCCHECK,
            CRC_ERR            => CRC_ERR
        );

    UUT_data_seq_check: entity work.data_seq_check
        port map (
            RST_N                  => RST_N,
            CLK                    => CLK,
            DATA_DCCHECK           => DATA_DCCHECK,
            SEQ_NUM_DCCHECK        => SEQ_NUM_DCCHECK,
            REC_POLARITY_FLG       => REC_POLARITY_FLG,
            END_FRAME_DCCHECK         => END_FRAME_DCCHECK,
            TYPE_FRAME_DCCHECK     => TYPE_FRAME_DCCHECK,
            NEW_WORD_DCCHECK       => NEW_WORD_DCCHECK,
            DATA_DSCHECK      => DATA_DSCHECK,
            NEW_WORD_DSCHECK       => NEW_WORD_DSCHECK,
            END_FRAME_DSCHECK         => END_FRAME_DSCHECK,
            SEQ_NUM_ERR            => SEQ_NUM_ERR,
            FIFO_FULL              => FIFO_FULL
        );

end Behavioral;
