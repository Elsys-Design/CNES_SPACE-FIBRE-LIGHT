----------------------------------------------------------------------------
-- Author(s) : Y. DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 24/02/2025
--
-- Description : This module checks the validity of the SEQ_num
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;



entity demux_rx is
  port (
    RST_N                  : in  std_logic; --! Global reset
    CLK                    : in  std_logic; --! Global Clock
    -- Ctrl signal
    ENABLE_SPY             : in std_logic;  --! Enable Spy read command
    -- Data-Link interface
    FIFO_RX_RD_EN_DL       : in  std_logic; --! Flag to read data in FIFO RX from Data-Link
		-- SPY interface
    FIFO_RX_RD_EN_SPY      : in  std_logic; --! Flag to read data in FIFO RX from Spy
    -- Phy Plus Lane interface
    FIFO_RX_RD_EN_DEMUX    : out std_logic  --! Flag to read data in FIFO RX to PPL
  );
end demux_rx;

architecture rtl of demux_rx is
---------------------------------------------------------
-----                  Declaration signals          -----
---------------------------------------------------------
begin

---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
---------------------------------------------------------
-- Process: p_mux
-- Description: Multiplex Injector and data_link signals
---------------------------------------------------------
p_mux: process(CLK, RST_N)
begin
	if RST_N = '0' then
	  FIFO_RX_RD_EN_DEMUX             <= '0';
	elsif rising_edge(CLK) then
    if ENABLE_SPY ='1' then
      FIFO_RX_RD_EN_DEMUX           <= FIFO_RX_RD_EN_SPY;
    else
      FIFO_RX_RD_EN_DEMUX           <= FIFO_RX_RD_EN_DL;
	  end if;
	end if;
end process p_mux;

end architecture rtl;