`include "B_IBUFDSE3_defines.vh"

reg [`IBUFDSE3_DATA_SZ-1:0] ATTR [0:`IBUFDSE3_ADDR_N-1];
reg [`IBUFDSE3__DIFF_TERM_SZ:1] DIFF_TERM_REG = DIFF_TERM;
reg [`IBUFDSE3__DQS_BIAS_SZ:1] DQS_BIAS_REG = DQS_BIAS;
reg [`IBUFDSE3__IBUF_LOW_PWR_SZ:1] IBUF_LOW_PWR_REG = IBUF_LOW_PWR;
reg [`IBUFDSE3__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IBUFDSE3__SIM_DEVICE_SZ:1] SIM_DEVICE_REG = SIM_DEVICE;
reg [`IBUFDSE3__SIM_INPUT_BUFFER_OFFSET_SZ-1:0] SIM_INPUT_BUFFER_OFFSET_REG = SIM_INPUT_BUFFER_OFFSET;
reg [`IBUFDSE3__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IBUFDSE3__DIFF_TERM] = DIFF_TERM;
  ATTR[`IBUFDSE3__DQS_BIAS] = DQS_BIAS;
  ATTR[`IBUFDSE3__IBUF_LOW_PWR] = IBUF_LOW_PWR;
  ATTR[`IBUFDSE3__IOSTANDARD] = IOSTANDARD;
  ATTR[`IBUFDSE3__SIM_DEVICE] = SIM_DEVICE;
  ATTR[`IBUFDSE3__SIM_INPUT_BUFFER_OFFSET] = SIM_INPUT_BUFFER_OFFSET;
  ATTR[`IBUFDSE3__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  DIFF_TERM_REG = ATTR[`IBUFDSE3__DIFF_TERM];
  DQS_BIAS_REG = ATTR[`IBUFDSE3__DQS_BIAS];
  IBUF_LOW_PWR_REG = ATTR[`IBUFDSE3__IBUF_LOW_PWR];
  IOSTANDARD_REG = ATTR[`IBUFDSE3__IOSTANDARD];
  SIM_DEVICE_REG = ATTR[`IBUFDSE3__SIM_DEVICE];
  SIM_INPUT_BUFFER_OFFSET_REG = ATTR[`IBUFDSE3__SIM_INPUT_BUFFER_OFFSET];
  USE_IBUFDISABLE_REG = ATTR[`IBUFDSE3__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IBUFDSE3_ADDR_SZ-1:0] addr;
  input  [`IBUFDSE3_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IBUFDSE3_DATA_SZ-1:0] read_attr;
  input  [`IBUFDSE3_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
