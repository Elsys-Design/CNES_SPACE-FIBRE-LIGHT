-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 22/07/2025
--
-- Description : This module detect the control words in the data flow
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_lane_ctrl_word_detect is
  port (
    RST_N                            : in  std_logic;                                          --! global reset
    CLK                              : in  std_logic;                                          --! Clock generated by HSSL IP
    -- ppl_64_lane_init_fsm (PLIF) interface
    NO_SIGNAL_PLCWD                  : out std_logic;                                          --! Flag no signal are received
    RX_NEW_WORD_PLCWD                : out std_logic_vector(1 downto 0);                       --! Flag new word has been received
    DETECTED_INIT1_PLCWD             : out std_logic_vector(1 downto 0);                       --! Flag INIT1 control word rxed
    DETECTED_INIT2_PLCWD             : out std_logic_vector(1 downto 0);                       --! Flag INIT2 control word rxed
    DETECTED_INIT3_PLCWD             : out std_logic_vector(1 downto 0);                       --! Flag INIT3 control word rxed
    DETECTED_INV_INIT1_PLCWD         : out std_logic_vector(1 downto 0);                       --! Flag INV_INIT1 control word rxed
    DETECTED_INV_INIT2_PLCWD         : out std_logic_vector(1 downto 0);                       --! Flag INV_INIT2 control word rxed
    DETECTED_RXERR_WORD_PLCWD        : out std_logic_vector(1 downto 0);                       --! Flag RXERR detected
    DETECTED_LOSS_SIGNAL_PLCWD       : out std_logic_vector(1 downto 0);                       --! Flag LOSS_SIGNAL detected
    DETECTED_STANDBY_PLCWD           : out std_logic_vector(1 downto 0);                       --! Flag STANDBY detected
    COMMA_K287_RXED_PLCWD            : out std_logic_vector(1 downto 0);                       --! Flag Comma K28.7 has been received
    CAPABILITY_PLCWD                 : out std_logic_vector(15 downto 0);                      --! Capability from INIT3 control word (31 downto 24) and (63 downto 56)
    SEND_RXERR_PLIF                  : in  std_logic_vector(1 downto 0);                       --! Flag send RXERR control word to Data-Link layer when FSM leave ACTIVE_ST
    NO_SIGNAL_DETECTION_ENABLED_PLIF : in  std_logic;                                          --! Flag to enable the no signal function
    ENABLE_TRANSM_DATA_PLIF          : in  std_logic_vector(1 downto 0);                       --! Flag to enable the transmision of data
    -- ppl_64_parallel_looback (PLPL) interface
    DATA_RX_PLPL                     : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! 64-bit data from ppl_64_parallel_looback
    VALID_K_CHARAC_PLPL               : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! 8-bit valid K character flags from ppl_64_parallel_looback
    DATA_RDY_PLPL                    : in  std_logic;                                          --! Data valid flag from ppl_64_parallel_looback
    -- DATA-LINK interface
    DATA_RX_PLCWD                    : out std_logic_vector(C_DATA_LENGTH-1 downto 0);          --! 64-bit data to Data-link layer
    VALID_K_CHARAC_PLCWD              : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0);  --! 8-bit valid K character flags to Data-link layer
    DATA_RDY_PLCWD                   : out std_logic_vector(1 downto 0)                         --! Data valid flag to Data-link layer
  );
end ppl_64_lane_ctrl_word_detect;

architecture rtl of ppl_64_lane_ctrl_word_detect is
---------------------------------------------------------
-----                  Signal declaration           -----
---------------------------------------------------------
signal enable_transm_data_r  : std_logic_vector(1 downto 0);
signal enable_transm_data_rr : std_logic_vector(1 downto 0);

-- First word signals
signal rx_new_word_fw           : std_logic;
signal detected_init1_fw        : std_logic;
signal detected_init2_fw        : std_logic;
signal detected_init3_fw        : std_logic;
signal detected_inv_init1_fw    : std_logic;
signal detected_inv_init2_fw    : std_logic;
signal comma_k287_rxed_fw       : std_logic;
signal detected_loss_signal_fw  : std_logic;
signal detected_standby_fw      : std_logic;
signal data_rx_dl_fw            : std_logic_vector(31 downto 0);
signal valid_k_charac_dl_fw     : std_logic_vector(3 downto 0);
signal data_rdy_dl_fw           : std_logic;
signal detected_rxerr_word_fw   : std_logic;
signal capability_fw            : std_logic_vector(7 downto 0);
-- Second word signals
signal rx_new_word_sw           : std_logic;
signal detected_init1_sw        : std_logic;
signal detected_init2_sw        : std_logic;
signal detected_init3_sw        : std_logic;
signal detected_inv_init1_sw    : std_logic;
signal detected_inv_init2_sw    : std_logic;
signal comma_k287_rxed_sw       : std_logic;
signal detected_loss_signal_sw  : std_logic;
signal detected_standby_sw      : std_logic;
signal data_rx_dl_sw            : std_logic_vector(31 downto 0);
signal valid_k_charac_dl_sw     : std_logic_vector(3 downto 0);
signal data_rdy_dl_sw           : std_logic;
signal detected_rxerr_word_sw   : std_logic;
signal capability_sw            : std_logic_vector(7 downto 0);


begin
---------------------------------------------------------
-----                  Assignment                   -----
---------------------------------------------------------
-- Outputs
DATA_RX_PLCWD              <= data_rx_dl_sw           & data_rx_dl_fw;
VALID_K_CHARAC_PLCWD        <= valid_k_charac_dl_sw    & valid_k_charac_dl_fw;
DATA_RDY_PLCWD             <= data_rdy_dl_sw          & data_rdy_dl_fw;
RX_NEW_WORD_PLCWD          <= rx_new_word_sw          & rx_new_word_fw;
DETECTED_INIT1_PLCWD       <= detected_init1_sw       & detected_init1_fw;
DETECTED_INIT2_PLCWD       <= detected_init2_sw       & detected_init2_fw;
DETECTED_INIT3_PLCWD       <= detected_init3_sw       & detected_init3_fw;
DETECTED_INV_INIT1_PLCWD   <= detected_inv_init1_sw   & detected_inv_init1_fw;
DETECTED_INV_INIT2_PLCWD   <= detected_inv_init2_sw   & detected_inv_init2_fw;
DETECTED_RXERR_WORD_PLCWD  <= detected_rxerr_word_sw  & detected_rxerr_word_fw;
DETECTED_LOSS_SIGNAL_PLCWD <= detected_loss_signal_sw & detected_loss_signal_fw;
DETECTED_STANDBY_PLCWD     <= detected_standby_sw     & detected_standby_fw;
COMMA_K287_RXED_PLCWD      <= comma_k287_rxed_sw      & comma_k287_rxed_fw;
CAPABILITY_PLCWD           <= capability_sw           & capability_fw;
---------------------------------------------------------
-----                     Process                   -----
---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_first_ctrl_word_detection
  -- Description: Detection of the control words for the first word.
  ---------------------------------------------------------
  p_first_ctrl_word_detection : process(CLK, RST_N)
  begin
    if RST_N = '0' then
      rx_new_word_fw           <= '0';
      detected_init1_fw        <= '0';
      detected_init2_fw        <= '0';
      detected_init3_fw        <= '0';
      detected_inv_init1_fw    <= '0';
      detected_inv_init2_fw    <= '0';
      comma_k287_rxed_fw       <= '0';
      detected_loss_signal_fw  <= '0';
      detected_standby_fw      <= '0';
      data_rx_dl_fw            <= (others => '0');
      valid_k_charac_dl_fw     <= (others => '0');
      data_rdy_dl_fw           <= '0';
      detected_rxerr_word_fw   <= '0';
      capability_fw            <= (others => '0');
    elsif rising_edge(CLK) then
      -- reset flags
      rx_new_word_fw          <= '0';
      detected_init1_fw       <= '0';
      detected_init2_fw       <= '0';
      detected_init3_fw       <= '0';
      detected_inv_init1_fw   <= '0';
      detected_inv_init2_fw   <= '0';
      comma_k287_rxed_fw      <= '0';
      detected_loss_signal_fw <= '0';
      detected_standby_fw     <= '0';
      capability_fw            <= (others => '0');
      data_rdy_dl_fw          <= '0';
      data_rx_dl_fw           <= (others => '0');
      valid_k_charac_dl_fw    <= (others => '0');
      detected_rxerr_word_fw  <= '0';
      -- Control word identification
      if DATA_RDY_PLPL = '1' then
        -- INIT 1
        if DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_INIT1_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_init1_fw   <= '1';
          rx_new_word_fw      <= '1';
        -- INIT 2
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_INIT2_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_init2_fw   <= '1';
          rx_new_word_fw      <= '1';
        -- INIT 3
        elsif DATA_RX_PLPL(23 downto 0) = C_INIT3_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_init3_fw   <= '1';
          rx_new_word_fw      <= '1';
          capability_fw       <= DATA_RX_PLPL(31 downto 24);
        -- iINIT 1
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_I_INIT1_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_inv_init1_fw <= '1';
          rx_new_word_fw        <= '1';
        -- iINIT 2
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_I_INIT2_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_inv_init2_fw <= '1';
          rx_new_word_fw        <= '1';
        -- LOST SIGNAL
        elsif DATA_RX_PLPL(23 downto 0) = C_LOST_SIG_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_loss_signal_fw <= '1';
          comma_k287_rxed_fw      <= '1';
          rx_new_word_fw          <= '1';
        -- STANDBY
        elsif DATA_RX_PLPL(23 downto 0) = C_STANDBY_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          detected_standby_fw    <= '1';
          comma_k287_rxed_fw     <= '1';
          rx_new_word_fw         <= '1';
        -- SEND RXERR
        elsif SEND_RXERR_PLIF(0) = '1' then
          data_rx_dl_fw        <= C_RXERR_WORD;
          valid_k_charac_dl_fw <= x"1";
          data_rdy_dl_fw       <= '1';
        -- Transmit DATA
        elsif enable_transm_data_rr(0) = '1' and not((DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_IDLE_WORD or DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_SKIP_WORD) and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1") then
          data_rx_dl_fw        <= DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0);
          valid_k_charac_dl_fw <= VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0);
          data_rdy_dl_fw       <= DATA_RDY_PLPL;
          rx_new_word_fw       <= '1';
          if DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_RXERR_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
            detected_rxerr_word_fw <= '1';
          end if;
        -- SKIP or IDLE
        elsif (DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_IDLE_WORD or DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_SKIP_WORD) and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
          comma_k287_rxed_fw   <= '1';
          rx_new_word_fw       <= '1';
        else
          rx_new_word_fw       <= '1';
          if DATA_RX_PLPL(C_DATA_LENGTH/2-1 downto 0) = C_RXERR_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH/2-1 downto 0) = x"1" then
            detected_rxerr_word_fw <= '1';
          end if;
        end if;
      end if;
    end if;
  end process p_first_ctrl_word_detection;
  ---------------------------------------------------------
  --! Process: p_second_ctrl_word_detection
  --! Description: Detection of the control words for the second word.
  ---------------------------------------------------------
  p_second_ctrl_word_detection : process(CLK, RST_N)
  begin
    if RST_N = '0' then
      rx_new_word_sw           <= '0';
      detected_init1_sw        <= '0';
      detected_init2_sw        <= '0';
      detected_init3_sw        <= '0';
      detected_inv_init1_sw    <= '0';
      detected_inv_init2_sw    <= '0';
      comma_k287_rxed_sw       <= '0';
      detected_loss_signal_sw  <= '0';
      detected_standby_sw      <= '0';
      data_rx_dl_sw            <= (others => '0');
      valid_k_charac_dl_sw     <= (others => '0');
      data_rdy_dl_sw           <= '0';
      detected_rxerr_word_sw   <= '0';
      capability_sw            <= (others => '0');
    elsif rising_edge(CLK) then
      -- reset flags
      rx_new_word_sw          <= '0';
      detected_init1_sw       <= '0';
      detected_init2_sw       <= '0';
      detected_init3_sw       <= '0';
      detected_inv_init1_sw   <= '0';
      detected_inv_init2_sw   <= '0';
      comma_k287_rxed_sw      <= '0';
      detected_loss_signal_sw <= '0';
      detected_standby_sw     <= '0';
      capability_sw           <= (others => '0');
      data_rdy_dl_sw          <= '0';
      data_rx_dl_sw           <= (others => '0');
      valid_k_charac_dl_sw    <= (others => '0');
      detected_rxerr_word_sw  <= '0';
      -- Control word identification
      if DATA_RDY_PLPL = '1' then
        -- INIT 1
        if DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_INIT1_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_init1_sw   <= '1';
          rx_new_word_sw      <= '1';
        -- INIT 2
        elsif DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_INIT2_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_init2_sw   <= '1';
          rx_new_word_sw      <= '1';
        -- INIT 3
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2+23 downto C_DATA_LENGTH/2) = C_INIT3_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_init3_sw   <= '1';
          rx_new_word_sw      <= '1';
          capability_sw       <= DATA_RX_PLPL(63 downto 56);
        -- iINIT 1
        elsif DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_I_INIT1_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_inv_init1_sw <= '1';
          rx_new_word_sw        <= '1';
        -- iINIT 2
        elsif DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_I_INIT2_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_inv_init2_sw <= '1';
          rx_new_word_sw        <= '1';
        -- LOST SIGNAL
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2+23 downto C_DATA_LENGTH/2) = C_LOST_SIG_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_loss_signal_sw <= '1';
          comma_k287_rxed_sw      <= '1';
          rx_new_word_sw          <= '1';
        -- STANDBY
        elsif DATA_RX_PLPL(C_DATA_LENGTH/2+23 downto C_DATA_LENGTH/2) = C_STANDBY_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          detected_standby_sw  <= '1';
          comma_k287_rxed_sw   <= '1';
          rx_new_word_sw       <= '1';
        -- SEND RXERR
        elsif SEND_RXERR_PLIF(1) = '1' then
          data_rx_dl_sw        <= C_RXERR_WORD;
          valid_k_charac_dl_sw <= x"1";
          data_rdy_dl_sw       <= '1';
        -- Transmit DATA
        elsif enable_transm_data_rr(1) = '1' and not((DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_IDLE_WORD or DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_SKIP_WORD) and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1") then
          data_rx_dl_sw        <= DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2);
          valid_k_charac_dl_sw <= VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2);
          data_rdy_dl_sw       <= DATA_RDY_PLPL;
          rx_new_word_sw       <= '1';
          if DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_RXERR_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
            detected_rxerr_word_sw <= '1';
          end if;
        -- SKIP or IDLE
        elsif (DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_IDLE_WORD or DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_SKIP_WORD) and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
          comma_k287_rxed_sw   <= '1';
          rx_new_word_sw       <= '1';
        else
          rx_new_word_sw       <= '1';
          if DATA_RX_PLPL(C_DATA_LENGTH-1 downto C_DATA_LENGTH/2) = C_RXERR_WORD and VALID_K_CHARAC_PLPL(C_BYTE_BY_WORD_LENGTH-1 downto C_BYTE_BY_WORD_LENGTH/2) = x"1" then
            detected_rxerr_word_sw <= '1';
          end if;
        end if;
      end if;
    end if;
  end process p_second_ctrl_word_detection;
  ---------------------------------------------------------
  -- Process: p_no_signal_detection
  -- Description: No signal detection.
  ---------------------------------------------------------
  p_no_signal_detection : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      NO_SIGNAL_PLCWD   <= '0';
    elsif rising_edge(CLK) then
      if NO_SIGNAL_DETECTION_ENABLED_PLIF = '1' then
        NO_SIGNAL_PLCWD   <= '1';
      else
        NO_SIGNAL_PLCWD   <= '0';
      end if;
    end if;
  end process p_no_signal_detection;

  ---------------------------------------------------------
  -- Process: p_enable_transm_data
  -- Description: ENABLE_TRANSM_DATA_PLIF delayed
  ---------------------------------------------------------
  p_enable_transm_data : process(CLK,RST_N)
  begin
    if RST_N = '0' then
      enable_transm_data_r     <= "00";
      enable_transm_data_rr    <= "00";
    elsif rising_edge(CLK) then
      enable_transm_data_r  <= ENABLE_TRANSM_DATA_PLIF;
      enable_transm_data_rr <= enable_transm_data_r;
    end if;
  end process p_enable_transm_data;
end architecture rtl;