-----------------------------------------------------------------------------------
-- #                          Copyright CNES 2025                                 #
-- #                                                                              #
-- # This source describes Open Hardware and is licensed under the CERN-OHL-W v2. #
-- #                                                                              #
-- # You may redistribute and modify this documentation and make products         #
-- # using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).     #
-- #                                                                              #
-- # This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED             #
-- # WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY                 #
-- # AND FITNESS FOR A PARTICULAR PURPOSE.                                        #
-- #                                                                              #
-- # Please see the CERN-OHL-W v2 for applicable conditions.                      #
-----------------------------------------------------------------------------------
----------------------------------------------------------------------------
-- Author(s) : Y.DAURIAC
--
-- Project : IP SpaceFibreLight
--
-- Creation date : 07/07/2025
--
-- Description : This module implements the skip insertion word function
----------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library phy_plus_lane_64_lib;
   use phy_plus_lane_64_lib.pkg_phy_plus_lane_64b.all;

entity ppl_64_skip_insertion is
   port (
      RST_N                   : in  std_logic;                                          --! Global reset (Active low)
      CLK                     : in  std_logic;                                          --! Clock generated by HSSL IP
      -- ppl_64_lane_ctrl_word_insert (PLCWI) Interface
      NEW_DATA_PLCWI          : in  std_logic;                                          --! New data Flag
      DATA_TX_PLCWI           : in  std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit receive from DATA_LINK layer
      VALID_K_CHARAC_PLCWI    : in  std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character from DATA-LINK layer
      WAIT_SEND_DATA_PLSI      : out std_logic;                                          --! Flag to indicates that the lane_ctrl_word_insert send a SKIP control word
      -- HSSL Interface
      DATA_TX_PSI             : out std_logic_vector(C_DATA_LENGTH-1 downto 0);         --! Data 64-bit send to manufacturer IP
      VALID_K_CHARAC_PSI      : out std_logic_vector(C_BYTE_BY_WORD_LENGTH-1 downto 0); --! Flags indicates which byte is a K character
      -- ppl_64_lane_init_fsm
      ENABLE_TRANSM_DATA_PLIF_PLIF : in  std_logic                                           --! Flag to enable to send data
   );
end ppl_64_skip_insertion;

architecture rtl of ppl_64_skip_insertion is
  ---------------------------------------------------------
  -----                   Type declaration            -----
  ----------------------------------------------------------
  type state_type is (TX_INIT_ST,
                      TX_DATA_1_ST,
                      TX_DATA_2_ST,
                      TX_SKIP_1_ST,
                      TX_SKIP_2_ST
                      );
  ---------------------------------------------------------
  -----                  Signal declaration           -----
  ---------------------------------------------------------
  signal data_2    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0);
  signal data_1    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0);
  signal data_0    : std_logic_vector(C_DATA_LENGTH/2-1 downto 0);

  signal k_char_2  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0);
  signal k_char_1  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0);
  signal k_char_0  : std_logic_vector(C_BYTE_BY_WORD_LENGTH/2-1 downto 0);

  signal state     : state_type;
  signal state_cnt : unsigned(13-1 downto 0);
begin
  ---------------------------------------------------------
  -----                     Assignement               -----
  ---------------------------------------------------------
  data_2   <= DATA_TX_PLCWI(C_DATA_LENGTH-1   downto C_DATA_LENGTH/2);
  data_1   <= DATA_TX_PLCWI(C_DATA_LENGTH/2-1 downto 0);
  k_char_2 <= VALID_K_CHARAC_PLCWI(C_BYTE_BY_WORD_LENGTH-1   downto C_BYTE_BY_WORD_LENGTH/2);
  k_char_1 <= VALID_K_CHARAC_PLCWI(C_BYTE_BY_WORD_LENGTH/2-1 downto 0);
  ---------------------------------------------------------
  -----                     Process                   -----
  ---------------------------------------------------------
  ---------------------------------------------------------
  -- Process: p_rx_sync_fsm_transition
  -- Description: Insert a skip word in the data flow every
  --              5000 words
  ---------------------------------------------------------
  p_skip_insertion: process(CLK,RST_N)
  begin
    if RST_N = '0' then
      state              <= TX_INIT_ST;
      state_cnt          <= (others => '0');
      data_0             <= (others => '0');
      k_char_0           <= (others => '0');
      DATA_TX_PSI        <= (others => '0');
      VALID_K_CHARAC_PSI <= (others => '0');
      WAIT_SEND_DATA_PLSI <= '0';
    elsif rising_edge(CLK) then
      data_0   <= data_2;
      k_char_0 <= k_char_2;
      case state is
        when TX_INIT_ST =>
                          DATA_TX_PSI        <= DATA_TX_PLCWI;
                          VALID_K_CHARAC_PSI <= VALID_K_CHARAC_PLCWI;
                          WAIT_SEND_DATA_PLSI <= '0';
                          state_cnt          <= (others => '0');
                          if ENABLE_TRANSM_DATA_PLIF_PLIF = '1' then -- When the lane_init_fsm is in ACTIVE_ST
                             state           <= TX_DATA_1_ST;
                          end if;

        when TX_DATA_1_ST =>
                          VALID_K_CHARAC_PSI <= k_char_2 & k_char_1;
                          DATA_TX_PSI        <= data_2 & data_1;
                          state_cnt          <= state_cnt + 2;
                          if ENABLE_TRANSM_DATA_PLIF_PLIF = '0' then -- When the lane_init_fsm is in ACTIVE_ST
                             state    <= TX_INIT_ST;
                          elsif state_cnt >= C_5000_WORDS then
                            state_cnt <= (others => '0');
                            state     <= TX_SKIP_1_ST;
                          end if;

        when TX_SKIP_1_ST =>
                          VALID_K_CHARAC_PSI <= k_char_1 & x"1";
                          DATA_TX_PSI        <= data_1 & C_SKIP_WORD;
                          state_cnt          <= state_cnt + 1;
                          state              <= TX_DATA_2_ST;

        when TX_DATA_2_ST =>
                          VALID_K_CHARAC_PSI    <= k_char_1 & k_char_0;
                          DATA_TX_PSI           <= data_1 & data_0;
                          state_cnt             <= state_cnt + 2;
                          if ENABLE_TRANSM_DATA_PLIF_PLIF = '0' then -- When the lane_init_fsm is in ACTIVE_ST
                             state              <= TX_INIT_ST;
                          elsif state_cnt >= C_5000_WORDS-1 then
                            state_cnt           <= (others => '0');
                            state               <= TX_SKIP_2_ST;
                            WAIT_SEND_DATA_PLSI  <= '1';
                          end if;

        when TX_SKIP_2_ST =>
                          VALID_K_CHARAC_PSI <= x"1" & k_char_0;
                          DATA_TX_PSI        <= C_SKIP_WORD & data_0;
                          state_cnt          <= (others => '0');
                          state              <= TX_DATA_1_ST;
                          WAIT_SEND_DATA_PLSI <= '0';

        when others =>
                          DATA_TX_PSI        <= DATA_TX_PLCWI;
                          VALID_K_CHARAC_PSI <= VALID_K_CHARAC_PLCWI;
                          WAIT_SEND_DATA_PLSI <= '0';
                          state_cnt          <= (others => '0');

      end case;
    end if;
  end process p_skip_insertion;

end architecture rtl;
