// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_BUFGCE_DIV_DEFINES_VH
`else
`define B_BUFGCE_DIV_DEFINES_VH

// Look-up table parameters
//

`define BUFGCE_DIV_ADDR_N  8
`define BUFGCE_DIV_ADDR_SZ 32
`define BUFGCE_DIV_DATA_SZ 144

// Attribute addresses
//

`define BUFGCE_DIV__BUFGCE_DIVIDE    32'h00000000
`define BUFGCE_DIV__BUFGCE_DIVIDE_SZ 32

`define BUFGCE_DIV__CE_TYPE    32'h00000001
`define BUFGCE_DIV__CE_TYPE_SZ 64

`define BUFGCE_DIV__HARDSYNC_CLR    32'h00000002
`define BUFGCE_DIV__HARDSYNC_CLR_SZ 40

`define BUFGCE_DIV__IS_CE_INVERTED    32'h00000003
`define BUFGCE_DIV__IS_CE_INVERTED_SZ 1

`define BUFGCE_DIV__IS_CLR_INVERTED    32'h00000004
`define BUFGCE_DIV__IS_CLR_INVERTED_SZ 1

`define BUFGCE_DIV__IS_I_INVERTED    32'h00000005
`define BUFGCE_DIV__IS_I_INVERTED_SZ 1

`define BUFGCE_DIV__SIM_DEVICE    32'h00000006
`define BUFGCE_DIV__SIM_DEVICE_SZ 144

`define BUFGCE_DIV__STARTUP_SYNC    32'h00000007
`define BUFGCE_DIV__STARTUP_SYNC_SZ 40

`endif  // B_BUFGCE_DIV_DEFINES_VH
