// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IOBUFDS_DCIEN_DEFINES_VH
`else
`define B_IOBUFDS_DCIEN_DEFINES_VH

// Look-up table parameters
//

`define IOBUFDS_DCIEN_ADDR_N  7
`define IOBUFDS_DCIEN_ADDR_SZ 32
`define IOBUFDS_DCIEN_DATA_SZ 144

// Attribute addresses
//

`define IOBUFDS_DCIEN__DIFF_TERM    32'h00000000
`define IOBUFDS_DCIEN__DIFF_TERM_SZ 40

`define IOBUFDS_DCIEN__DQS_BIAS    32'h00000001
`define IOBUFDS_DCIEN__DQS_BIAS_SZ 40

`define IOBUFDS_DCIEN__IBUF_LOW_PWR    32'h00000002
`define IOBUFDS_DCIEN__IBUF_LOW_PWR_SZ 40

`define IOBUFDS_DCIEN__IOSTANDARD    32'h00000003
`define IOBUFDS_DCIEN__IOSTANDARD_SZ 56

`define IOBUFDS_DCIEN__SIM_DEVICE    32'h00000004
`define IOBUFDS_DCIEN__SIM_DEVICE_SZ 144

`define IOBUFDS_DCIEN__SLEW    32'h00000005
`define IOBUFDS_DCIEN__SLEW_SZ 48

`define IOBUFDS_DCIEN__USE_IBUFDISABLE    32'h00000006
`define IOBUFDS_DCIEN__USE_IBUFDISABLE_SZ 72

`endif  // B_IOBUFDS_DCIEN_DEFINES_VH