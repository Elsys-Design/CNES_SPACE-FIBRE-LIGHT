// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_MMCME3_ADV_DEFINES_VH
`else
`define B_MMCME3_ADV_DEFINES_VH

// Look-up table parameters
//

`define MMCME3_ADV_ADDR_N  57
`define MMCME3_ADV_ADDR_SZ 32
`define MMCME3_ADV_DATA_SZ 88

// Attribute addresses
//

`define MMCME3_ADV__BANDWIDTH    32'h00000000
`define MMCME3_ADV__BANDWIDTH_SZ 72

`define MMCME3_ADV__CLKFBOUT_MULT_F    32'h00000001
`define MMCME3_ADV__CLKFBOUT_MULT_F_SZ 64

`define MMCME3_ADV__CLKFBOUT_PHASE    32'h00000002
`define MMCME3_ADV__CLKFBOUT_PHASE_SZ 64

`define MMCME3_ADV__CLKFBOUT_USE_FINE_PS    32'h00000003
`define MMCME3_ADV__CLKFBOUT_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKIN1_PERIOD    32'h00000004
`define MMCME3_ADV__CLKIN1_PERIOD_SZ 64

`define MMCME3_ADV__CLKIN2_PERIOD    32'h00000005
`define MMCME3_ADV__CLKIN2_PERIOD_SZ 64

`define MMCME3_ADV__CLKIN_FREQ_MAX    32'h00000006
`define MMCME3_ADV__CLKIN_FREQ_MAX_SZ 64

`define MMCME3_ADV__CLKIN_FREQ_MIN    32'h00000007
`define MMCME3_ADV__CLKIN_FREQ_MIN_SZ 64

`define MMCME3_ADV__CLKOUT0_DIVIDE_F    32'h00000008
`define MMCME3_ADV__CLKOUT0_DIVIDE_F_SZ 64

`define MMCME3_ADV__CLKOUT0_DUTY_CYCLE    32'h00000009
`define MMCME3_ADV__CLKOUT0_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT0_PHASE    32'h0000000a
`define MMCME3_ADV__CLKOUT0_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT0_USE_FINE_PS    32'h0000000b
`define MMCME3_ADV__CLKOUT0_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT1_DIVIDE    32'h0000000c
`define MMCME3_ADV__CLKOUT1_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT1_DUTY_CYCLE    32'h0000000d
`define MMCME3_ADV__CLKOUT1_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT1_PHASE    32'h0000000e
`define MMCME3_ADV__CLKOUT1_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT1_USE_FINE_PS    32'h0000000f
`define MMCME3_ADV__CLKOUT1_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT2_DIVIDE    32'h00000010
`define MMCME3_ADV__CLKOUT2_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT2_DUTY_CYCLE    32'h00000011
`define MMCME3_ADV__CLKOUT2_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT2_PHASE    32'h00000012
`define MMCME3_ADV__CLKOUT2_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT2_USE_FINE_PS    32'h00000013
`define MMCME3_ADV__CLKOUT2_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT3_DIVIDE    32'h00000014
`define MMCME3_ADV__CLKOUT3_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT3_DUTY_CYCLE    32'h00000015
`define MMCME3_ADV__CLKOUT3_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT3_PHASE    32'h00000016
`define MMCME3_ADV__CLKOUT3_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT3_USE_FINE_PS    32'h00000017
`define MMCME3_ADV__CLKOUT3_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT4_CASCADE    32'h00000018
`define MMCME3_ADV__CLKOUT4_CASCADE_SZ 40

`define MMCME3_ADV__CLKOUT4_DIVIDE    32'h00000019
`define MMCME3_ADV__CLKOUT4_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT4_DUTY_CYCLE    32'h0000001a
`define MMCME3_ADV__CLKOUT4_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT4_PHASE    32'h0000001b
`define MMCME3_ADV__CLKOUT4_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT4_USE_FINE_PS    32'h0000001c
`define MMCME3_ADV__CLKOUT4_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT5_DIVIDE    32'h0000001d
`define MMCME3_ADV__CLKOUT5_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT5_DUTY_CYCLE    32'h0000001e
`define MMCME3_ADV__CLKOUT5_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT5_PHASE    32'h0000001f
`define MMCME3_ADV__CLKOUT5_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT5_USE_FINE_PS    32'h00000020
`define MMCME3_ADV__CLKOUT5_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKOUT6_DIVIDE    32'h00000021
`define MMCME3_ADV__CLKOUT6_DIVIDE_SZ 32

`define MMCME3_ADV__CLKOUT6_DUTY_CYCLE    32'h00000022
`define MMCME3_ADV__CLKOUT6_DUTY_CYCLE_SZ 64

`define MMCME3_ADV__CLKOUT6_PHASE    32'h00000023
`define MMCME3_ADV__CLKOUT6_PHASE_SZ 64

`define MMCME3_ADV__CLKOUT6_USE_FINE_PS    32'h00000024
`define MMCME3_ADV__CLKOUT6_USE_FINE_PS_SZ 40

`define MMCME3_ADV__CLKPFD_FREQ_MAX    32'h00000025
`define MMCME3_ADV__CLKPFD_FREQ_MAX_SZ 64

`define MMCME3_ADV__CLKPFD_FREQ_MIN    32'h00000026
`define MMCME3_ADV__CLKPFD_FREQ_MIN_SZ 64

`define MMCME3_ADV__COMPENSATION    32'h00000027
`define MMCME3_ADV__COMPENSATION_SZ 64

`define MMCME3_ADV__DIVCLK_DIVIDE    32'h00000028
`define MMCME3_ADV__DIVCLK_DIVIDE_SZ 32

`define MMCME3_ADV__IS_CLKFBIN_INVERTED    32'h00000029
`define MMCME3_ADV__IS_CLKFBIN_INVERTED_SZ 1

`define MMCME3_ADV__IS_CLKIN1_INVERTED    32'h0000002a
`define MMCME3_ADV__IS_CLKIN1_INVERTED_SZ 1

`define MMCME3_ADV__IS_CLKIN2_INVERTED    32'h0000002b
`define MMCME3_ADV__IS_CLKIN2_INVERTED_SZ 1

`define MMCME3_ADV__IS_CLKINSEL_INVERTED    32'h0000002c
`define MMCME3_ADV__IS_CLKINSEL_INVERTED_SZ 1

`define MMCME3_ADV__IS_PSEN_INVERTED    32'h0000002d
`define MMCME3_ADV__IS_PSEN_INVERTED_SZ 1

`define MMCME3_ADV__IS_PSINCDEC_INVERTED    32'h0000002e
`define MMCME3_ADV__IS_PSINCDEC_INVERTED_SZ 1

`define MMCME3_ADV__IS_PWRDWN_INVERTED    32'h0000002f
`define MMCME3_ADV__IS_PWRDWN_INVERTED_SZ 1

`define MMCME3_ADV__IS_RST_INVERTED    32'h00000030
`define MMCME3_ADV__IS_RST_INVERTED_SZ 1

`define MMCME3_ADV__REF_JITTER1    32'h00000031
`define MMCME3_ADV__REF_JITTER1_SZ 64

`define MMCME3_ADV__REF_JITTER2    32'h00000032
`define MMCME3_ADV__REF_JITTER2_SZ 64

`define MMCME3_ADV__SS_EN    32'h00000033
`define MMCME3_ADV__SS_EN_SZ 40

`define MMCME3_ADV__SS_MODE    32'h00000034
`define MMCME3_ADV__SS_MODE_SZ 88

`define MMCME3_ADV__SS_MOD_PERIOD    32'h00000035
`define MMCME3_ADV__SS_MOD_PERIOD_SZ 32

`define MMCME3_ADV__STARTUP_WAIT    32'h00000036
`define MMCME3_ADV__STARTUP_WAIT_SZ 40

`define MMCME3_ADV__VCOCLK_FREQ_MAX    32'h00000037
`define MMCME3_ADV__VCOCLK_FREQ_MAX_SZ 64

`define MMCME3_ADV__VCOCLK_FREQ_MIN    32'h00000038
`define MMCME3_ADV__VCOCLK_FREQ_MIN_SZ 64

`endif  // B_MMCME3_ADV_DEFINES_VH