// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_RAMB18E1_DEFINES_VH
`else
`define B_RAMB18E1_DEFINES_VH

// Look-up table parameters
//

`define RAMB18E1_ADDR_N  99
`define RAMB18E1_ADDR_SZ 32
`define RAMB18E1_DATA_SZ 256

// Attribute addresses
//

`define RAMB18E1__DOA_REG    32'h00000000
`define RAMB18E1__DOA_REG_SZ 32

`define RAMB18E1__DOB_REG    32'h00000001
`define RAMB18E1__DOB_REG_SZ 32

`define RAMB18E1__INITP_00    32'h00000002
`define RAMB18E1__INITP_00_SZ 256

`define RAMB18E1__INITP_01    32'h00000003
`define RAMB18E1__INITP_01_SZ 256

`define RAMB18E1__INITP_02    32'h00000004
`define RAMB18E1__INITP_02_SZ 256

`define RAMB18E1__INITP_03    32'h00000005
`define RAMB18E1__INITP_03_SZ 256

`define RAMB18E1__INITP_04    32'h00000006
`define RAMB18E1__INITP_04_SZ 256

`define RAMB18E1__INITP_05    32'h00000007
`define RAMB18E1__INITP_05_SZ 256

`define RAMB18E1__INITP_06    32'h00000008
`define RAMB18E1__INITP_06_SZ 256

`define RAMB18E1__INITP_07    32'h00000009
`define RAMB18E1__INITP_07_SZ 256

`define RAMB18E1__INIT_00    32'h0000000a
`define RAMB18E1__INIT_00_SZ 256

`define RAMB18E1__INIT_01    32'h0000000b
`define RAMB18E1__INIT_01_SZ 256

`define RAMB18E1__INIT_02    32'h0000000c
`define RAMB18E1__INIT_02_SZ 256

`define RAMB18E1__INIT_03    32'h0000000d
`define RAMB18E1__INIT_03_SZ 256

`define RAMB18E1__INIT_04    32'h0000000e
`define RAMB18E1__INIT_04_SZ 256

`define RAMB18E1__INIT_05    32'h0000000f
`define RAMB18E1__INIT_05_SZ 256

`define RAMB18E1__INIT_06    32'h00000010
`define RAMB18E1__INIT_06_SZ 256

`define RAMB18E1__INIT_07    32'h00000011
`define RAMB18E1__INIT_07_SZ 256

`define RAMB18E1__INIT_08    32'h00000012
`define RAMB18E1__INIT_08_SZ 256

`define RAMB18E1__INIT_09    32'h00000013
`define RAMB18E1__INIT_09_SZ 256

`define RAMB18E1__INIT_0A    32'h00000014
`define RAMB18E1__INIT_0A_SZ 256

`define RAMB18E1__INIT_0B    32'h00000015
`define RAMB18E1__INIT_0B_SZ 256

`define RAMB18E1__INIT_0C    32'h00000016
`define RAMB18E1__INIT_0C_SZ 256

`define RAMB18E1__INIT_0D    32'h00000017
`define RAMB18E1__INIT_0D_SZ 256

`define RAMB18E1__INIT_0E    32'h00000018
`define RAMB18E1__INIT_0E_SZ 256

`define RAMB18E1__INIT_0F    32'h00000019
`define RAMB18E1__INIT_0F_SZ 256

`define RAMB18E1__INIT_10    32'h0000001a
`define RAMB18E1__INIT_10_SZ 256

`define RAMB18E1__INIT_11    32'h0000001b
`define RAMB18E1__INIT_11_SZ 256

`define RAMB18E1__INIT_12    32'h0000001c
`define RAMB18E1__INIT_12_SZ 256

`define RAMB18E1__INIT_13    32'h0000001d
`define RAMB18E1__INIT_13_SZ 256

`define RAMB18E1__INIT_14    32'h0000001e
`define RAMB18E1__INIT_14_SZ 256

`define RAMB18E1__INIT_15    32'h0000001f
`define RAMB18E1__INIT_15_SZ 256

`define RAMB18E1__INIT_16    32'h00000020
`define RAMB18E1__INIT_16_SZ 256

`define RAMB18E1__INIT_17    32'h00000021
`define RAMB18E1__INIT_17_SZ 256

`define RAMB18E1__INIT_18    32'h00000022
`define RAMB18E1__INIT_18_SZ 256

`define RAMB18E1__INIT_19    32'h00000023
`define RAMB18E1__INIT_19_SZ 256

`define RAMB18E1__INIT_1A    32'h00000024
`define RAMB18E1__INIT_1A_SZ 256

`define RAMB18E1__INIT_1B    32'h00000025
`define RAMB18E1__INIT_1B_SZ 256

`define RAMB18E1__INIT_1C    32'h00000026
`define RAMB18E1__INIT_1C_SZ 256

`define RAMB18E1__INIT_1D    32'h00000027
`define RAMB18E1__INIT_1D_SZ 256

`define RAMB18E1__INIT_1E    32'h00000028
`define RAMB18E1__INIT_1E_SZ 256

`define RAMB18E1__INIT_1F    32'h00000029
`define RAMB18E1__INIT_1F_SZ 256

`define RAMB18E1__INIT_20    32'h0000002a
`define RAMB18E1__INIT_20_SZ 256

`define RAMB18E1__INIT_21    32'h0000002b
`define RAMB18E1__INIT_21_SZ 256

`define RAMB18E1__INIT_22    32'h0000002c
`define RAMB18E1__INIT_22_SZ 256

`define RAMB18E1__INIT_23    32'h0000002d
`define RAMB18E1__INIT_23_SZ 256

`define RAMB18E1__INIT_24    32'h0000002e
`define RAMB18E1__INIT_24_SZ 256

`define RAMB18E1__INIT_25    32'h0000002f
`define RAMB18E1__INIT_25_SZ 256

`define RAMB18E1__INIT_26    32'h00000030
`define RAMB18E1__INIT_26_SZ 256

`define RAMB18E1__INIT_27    32'h00000031
`define RAMB18E1__INIT_27_SZ 256

`define RAMB18E1__INIT_28    32'h00000032
`define RAMB18E1__INIT_28_SZ 256

`define RAMB18E1__INIT_29    32'h00000033
`define RAMB18E1__INIT_29_SZ 256

`define RAMB18E1__INIT_2A    32'h00000034
`define RAMB18E1__INIT_2A_SZ 256

`define RAMB18E1__INIT_2B    32'h00000035
`define RAMB18E1__INIT_2B_SZ 256

`define RAMB18E1__INIT_2C    32'h00000036
`define RAMB18E1__INIT_2C_SZ 256

`define RAMB18E1__INIT_2D    32'h00000037
`define RAMB18E1__INIT_2D_SZ 256

`define RAMB18E1__INIT_2E    32'h00000038
`define RAMB18E1__INIT_2E_SZ 256

`define RAMB18E1__INIT_2F    32'h00000039
`define RAMB18E1__INIT_2F_SZ 256

`define RAMB18E1__INIT_30    32'h0000003a
`define RAMB18E1__INIT_30_SZ 256

`define RAMB18E1__INIT_31    32'h0000003b
`define RAMB18E1__INIT_31_SZ 256

`define RAMB18E1__INIT_32    32'h0000003c
`define RAMB18E1__INIT_32_SZ 256

`define RAMB18E1__INIT_33    32'h0000003d
`define RAMB18E1__INIT_33_SZ 256

`define RAMB18E1__INIT_34    32'h0000003e
`define RAMB18E1__INIT_34_SZ 256

`define RAMB18E1__INIT_35    32'h0000003f
`define RAMB18E1__INIT_35_SZ 256

`define RAMB18E1__INIT_36    32'h00000040
`define RAMB18E1__INIT_36_SZ 256

`define RAMB18E1__INIT_37    32'h00000041
`define RAMB18E1__INIT_37_SZ 256

`define RAMB18E1__INIT_38    32'h00000042
`define RAMB18E1__INIT_38_SZ 256

`define RAMB18E1__INIT_39    32'h00000043
`define RAMB18E1__INIT_39_SZ 256

`define RAMB18E1__INIT_3A    32'h00000044
`define RAMB18E1__INIT_3A_SZ 256

`define RAMB18E1__INIT_3B    32'h00000045
`define RAMB18E1__INIT_3B_SZ 256

`define RAMB18E1__INIT_3C    32'h00000046
`define RAMB18E1__INIT_3C_SZ 256

`define RAMB18E1__INIT_3D    32'h00000047
`define RAMB18E1__INIT_3D_SZ 256

`define RAMB18E1__INIT_3E    32'h00000048
`define RAMB18E1__INIT_3E_SZ 256

`define RAMB18E1__INIT_3F    32'h00000049
`define RAMB18E1__INIT_3F_SZ 256

`define RAMB18E1__INIT_A    32'h0000004a
`define RAMB18E1__INIT_A_SZ 18

`define RAMB18E1__INIT_B    32'h0000004b
`define RAMB18E1__INIT_B_SZ 18

`define RAMB18E1__INIT_FILE    32'h0000004c
`define RAMB18E1__INIT_FILE_SZ 32

`define RAMB18E1__IS_CLKARDCLK_INVERTED    32'h0000004d
`define RAMB18E1__IS_CLKARDCLK_INVERTED_SZ 1

`define RAMB18E1__IS_CLKBWRCLK_INVERTED    32'h0000004e
`define RAMB18E1__IS_CLKBWRCLK_INVERTED_SZ 1

`define RAMB18E1__IS_ENARDEN_INVERTED    32'h0000004f
`define RAMB18E1__IS_ENARDEN_INVERTED_SZ 1

`define RAMB18E1__IS_ENBWREN_INVERTED    32'h00000050
`define RAMB18E1__IS_ENBWREN_INVERTED_SZ 1

`define RAMB18E1__IS_RSTRAMARSTRAM_INVERTED    32'h00000051
`define RAMB18E1__IS_RSTRAMARSTRAM_INVERTED_SZ 1

`define RAMB18E1__IS_RSTRAMB_INVERTED    32'h00000052
`define RAMB18E1__IS_RSTRAMB_INVERTED_SZ 1

`define RAMB18E1__IS_RSTREGARSTREG_INVERTED    32'h00000053
`define RAMB18E1__IS_RSTREGARSTREG_INVERTED_SZ 1

`define RAMB18E1__IS_RSTREGB_INVERTED    32'h00000054
`define RAMB18E1__IS_RSTREGB_INVERTED_SZ 1

`define RAMB18E1__RAM_MODE    32'h00000055
`define RAMB18E1__RAM_MODE_SZ 24

`define RAMB18E1__RDADDR_COLLISION_HWCONFIG    32'h00000056
`define RAMB18E1__RDADDR_COLLISION_HWCONFIG_SZ 104

`define RAMB18E1__READ_WIDTH_A    32'h00000057
`define RAMB18E1__READ_WIDTH_A_SZ 32

`define RAMB18E1__READ_WIDTH_B    32'h00000058
`define RAMB18E1__READ_WIDTH_B_SZ 32

`define RAMB18E1__RSTREG_PRIORITY_A    32'h00000059
`define RAMB18E1__RSTREG_PRIORITY_A_SZ 48

`define RAMB18E1__RSTREG_PRIORITY_B    32'h0000005a
`define RAMB18E1__RSTREG_PRIORITY_B_SZ 48

`define RAMB18E1__SIM_COLLISION_CHECK    32'h0000005b
`define RAMB18E1__SIM_COLLISION_CHECK_SZ 120

`define RAMB18E1__SIM_DEVICE    32'h0000005c
`define RAMB18E1__SIM_DEVICE_SZ 56

`define RAMB18E1__SRVAL_A    32'h0000005d
`define RAMB18E1__SRVAL_A_SZ 18

`define RAMB18E1__SRVAL_B    32'h0000005e
`define RAMB18E1__SRVAL_B_SZ 18

`define RAMB18E1__WRITE_MODE_A    32'h0000005f
`define RAMB18E1__WRITE_MODE_A_SZ 88

`define RAMB18E1__WRITE_MODE_B    32'h00000060
`define RAMB18E1__WRITE_MODE_B_SZ 88

`define RAMB18E1__WRITE_WIDTH_A    32'h00000061
`define RAMB18E1__WRITE_WIDTH_A_SZ 32

`define RAMB18E1__WRITE_WIDTH_B    32'h00000062
`define RAMB18E1__WRITE_WIDTH_B_SZ 32

`endif  // B_RAMB18E1_DEFINES_VH