`include "B_IOBUFDS_ODDR_defines.vh"

reg [`IOBUFDS_ODDR_DATA_SZ-1:0] ATTR [0:`IOBUFDS_ODDR_ADDR_N-1];
reg [`IOBUFDS_ODDR__DIFF_TERM_SZ:1] DIFF_TERM_REG = DIFF_TERM;
reg [`IOBUFDS_ODDR__DQS_BIAS_SZ:1] DQS_BIAS_REG = DQS_BIAS;
reg [`IOBUFDS_ODDR__EN_OMUX_SZ:1] EN_OMUX_REG = EN_OMUX;
reg [`IOBUFDS_ODDR__IOSTANDARD_SZ:1] IOSTANDARD_REG = IOSTANDARD;
reg [`IOBUFDS_ODDR__SIM_INPUT_BUFFER_OFFSET_SZ-1:0] SIM_INPUT_BUFFER_OFFSET_REG = SIM_INPUT_BUFFER_OFFSET;
reg [`IOBUFDS_ODDR__USE_IBUFDISABLE_SZ:1] USE_IBUFDISABLE_REG = USE_IBUFDISABLE;

initial begin
  ATTR[`IOBUFDS_ODDR__DIFF_TERM] = DIFF_TERM;
  ATTR[`IOBUFDS_ODDR__DQS_BIAS] = DQS_BIAS;
  ATTR[`IOBUFDS_ODDR__EN_OMUX] = EN_OMUX;
  ATTR[`IOBUFDS_ODDR__IOSTANDARD] = IOSTANDARD;
  ATTR[`IOBUFDS_ODDR__SIM_INPUT_BUFFER_OFFSET] = SIM_INPUT_BUFFER_OFFSET;
  ATTR[`IOBUFDS_ODDR__USE_IBUFDISABLE] = USE_IBUFDISABLE;
end

always @(trig_attr) begin
  DIFF_TERM_REG = ATTR[`IOBUFDS_ODDR__DIFF_TERM];
  DQS_BIAS_REG = ATTR[`IOBUFDS_ODDR__DQS_BIAS];
  EN_OMUX_REG = ATTR[`IOBUFDS_ODDR__EN_OMUX];
  IOSTANDARD_REG = ATTR[`IOBUFDS_ODDR__IOSTANDARD];
  SIM_INPUT_BUFFER_OFFSET_REG = ATTR[`IOBUFDS_ODDR__SIM_INPUT_BUFFER_OFFSET];
  USE_IBUFDISABLE_REG = ATTR[`IOBUFDS_ODDR__USE_IBUFDISABLE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`IOBUFDS_ODDR_ADDR_SZ-1:0] addr;
  input  [`IOBUFDS_ODDR_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`IOBUFDS_ODDR_DATA_SZ-1:0] read_attr;
  input  [`IOBUFDS_ODDR_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
trig_attr = ~trig_attr;
  end
endtask
