// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_XPLL_DEFINES_VH
`else
`define B_XPLL_DEFINES_VH

// Look-up table parameters
//

`define XPLL_ADDR_N  52
`define XPLL_ADDR_SZ 32
`define XPLL_DATA_SZ 64

// Attribute addresses
//

`define XPLL__CLKFBOUT_MULT    32'h00000000
`define XPLL__CLKFBOUT_MULT_SZ 32

`define XPLL__CLKFBOUT_PHASE    32'h00000001
`define XPLL__CLKFBOUT_PHASE_SZ 64

`define XPLL__CLKIN_FREQ_MAX    32'h00000002
`define XPLL__CLKIN_FREQ_MAX_SZ 64

`define XPLL__CLKIN_FREQ_MIN    32'h00000003
`define XPLL__CLKIN_FREQ_MIN_SZ 64

`define XPLL__CLKIN_PERIOD    32'h00000004
`define XPLL__CLKIN_PERIOD_SZ 64

`define XPLL__CLKOUT0_DIVIDE    32'h00000005
`define XPLL__CLKOUT0_DIVIDE_SZ 32

`define XPLL__CLKOUT0_DUTY_CYCLE    32'h00000006
`define XPLL__CLKOUT0_DUTY_CYCLE_SZ 64

`define XPLL__CLKOUT0_PHASE    32'h00000007
`define XPLL__CLKOUT0_PHASE_SZ 64

`define XPLL__CLKOUT0_PHASE_CTRL    32'h00000008
`define XPLL__CLKOUT0_PHASE_CTRL_SZ 2

`define XPLL__CLKOUT1_DIVIDE    32'h00000009
`define XPLL__CLKOUT1_DIVIDE_SZ 32

`define XPLL__CLKOUT1_DUTY_CYCLE    32'h0000000a
`define XPLL__CLKOUT1_DUTY_CYCLE_SZ 64

`define XPLL__CLKOUT1_PHASE    32'h0000000b
`define XPLL__CLKOUT1_PHASE_SZ 64

`define XPLL__CLKOUT1_PHASE_CTRL    32'h0000000c
`define XPLL__CLKOUT1_PHASE_CTRL_SZ 2

`define XPLL__CLKOUT2_DIVIDE    32'h0000000d
`define XPLL__CLKOUT2_DIVIDE_SZ 32

`define XPLL__CLKOUT2_DUTY_CYCLE    32'h0000000e
`define XPLL__CLKOUT2_DUTY_CYCLE_SZ 64

`define XPLL__CLKOUT2_PHASE    32'h0000000f
`define XPLL__CLKOUT2_PHASE_SZ 64

`define XPLL__CLKOUT2_PHASE_CTRL    32'h00000010
`define XPLL__CLKOUT2_PHASE_CTRL_SZ 2

`define XPLL__CLKOUT3_DIVIDE    32'h00000011
`define XPLL__CLKOUT3_DIVIDE_SZ 32

`define XPLL__CLKOUT3_DUTY_CYCLE    32'h00000012
`define XPLL__CLKOUT3_DUTY_CYCLE_SZ 64

`define XPLL__CLKOUT3_PHASE    32'h00000013
`define XPLL__CLKOUT3_PHASE_SZ 64

`define XPLL__CLKOUT3_PHASE_CTRL    32'h00000014
`define XPLL__CLKOUT3_PHASE_CTRL_SZ 2

`define XPLL__CLKOUTPHY_CASCIN_EN    32'h00000015
`define XPLL__CLKOUTPHY_CASCIN_EN_SZ 1

`define XPLL__CLKOUTPHY_CASCOUT_EN    32'h00000016
`define XPLL__CLKOUTPHY_CASCOUT_EN_SZ 1

`define XPLL__CLKOUTPHY_DIVIDE    32'h00000017
`define XPLL__CLKOUTPHY_DIVIDE_SZ 40

`define XPLL__CLKPFD_FREQ_MAX    32'h00000018
`define XPLL__CLKPFD_FREQ_MAX_SZ 64

`define XPLL__CLKPFD_FREQ_MIN    32'h00000019
`define XPLL__CLKPFD_FREQ_MIN_SZ 64

`define XPLL__DESKEW2_MUXIN_SEL    32'h0000001a
`define XPLL__DESKEW2_MUXIN_SEL_SZ 1

`define XPLL__DESKEW_DELAY1    32'h0000001b
`define XPLL__DESKEW_DELAY1_SZ 32

`define XPLL__DESKEW_DELAY2    32'h0000001c
`define XPLL__DESKEW_DELAY2_SZ 32

`define XPLL__DESKEW_DELAY_EN1    32'h0000001d
`define XPLL__DESKEW_DELAY_EN1_SZ 40

`define XPLL__DESKEW_DELAY_EN2    32'h0000001e
`define XPLL__DESKEW_DELAY_EN2_SZ 40

`define XPLL__DESKEW_DELAY_PATH1    32'h0000001f
`define XPLL__DESKEW_DELAY_PATH1_SZ 40

`define XPLL__DESKEW_DELAY_PATH2    32'h00000020
`define XPLL__DESKEW_DELAY_PATH2_SZ 40

`define XPLL__DESKEW_MUXIN_SEL    32'h00000021
`define XPLL__DESKEW_MUXIN_SEL_SZ 1

`define XPLL__DIV4_CLKOUT012    32'h00000022
`define XPLL__DIV4_CLKOUT012_SZ 1

`define XPLL__DIV4_CLKOUT3    32'h00000023
`define XPLL__DIV4_CLKOUT3_SZ 1

`define XPLL__DIVCLK_DIVIDE    32'h00000024
`define XPLL__DIVCLK_DIVIDE_SZ 32

`define XPLL__IS_CLKFB1_DESKEW_INVERTED    32'h00000025
`define XPLL__IS_CLKFB1_DESKEW_INVERTED_SZ 1

`define XPLL__IS_CLKFB2_DESKEW_INVERTED    32'h00000026
`define XPLL__IS_CLKFB2_DESKEW_INVERTED_SZ 1

`define XPLL__IS_CLKIN1_DESKEW_INVERTED    32'h00000027
`define XPLL__IS_CLKIN1_DESKEW_INVERTED_SZ 1

`define XPLL__IS_CLKIN2_DESKEW_INVERTED    32'h00000028
`define XPLL__IS_CLKIN2_DESKEW_INVERTED_SZ 1

`define XPLL__IS_CLKIN_INVERTED    32'h00000029
`define XPLL__IS_CLKIN_INVERTED_SZ 1

`define XPLL__IS_PSEN_INVERTED    32'h0000002a
`define XPLL__IS_PSEN_INVERTED_SZ 1

`define XPLL__IS_PSINCDEC_INVERTED    32'h0000002b
`define XPLL__IS_PSINCDEC_INVERTED_SZ 1

`define XPLL__IS_PWRDWN_INVERTED    32'h0000002c
`define XPLL__IS_PWRDWN_INVERTED_SZ 1

`define XPLL__IS_RST_INVERTED    32'h0000002d
`define XPLL__IS_RST_INVERTED_SZ 1

`define XPLL__LOCK_WAIT    32'h0000002e
`define XPLL__LOCK_WAIT_SZ 40

`define XPLL__REF_JITTER    32'h0000002f
`define XPLL__REF_JITTER_SZ 64

`define XPLL__SIM_ADJ_CLK0_CASCADE    32'h00000030
`define XPLL__SIM_ADJ_CLK0_CASCADE_SZ 40

`define XPLL__VCOCLK_FREQ_MAX    32'h00000031
`define XPLL__VCOCLK_FREQ_MAX_SZ 64

`define XPLL__VCOCLK_FREQ_MIN    32'h00000032
`define XPLL__VCOCLK_FREQ_MIN_SZ 64

`define XPLL__XPLL_CONNECT_TO_NOCMC    32'h00000033
`define XPLL__XPLL_CONNECT_TO_NOCMC_SZ 32

`endif  // B_XPLL_DEFINES_VH