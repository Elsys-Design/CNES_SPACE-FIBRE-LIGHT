// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_URAM288_BASE_DEFINES_VH
`else
`define B_URAM288_BASE_DEFINES_VH

// Look-up table parameters
//

`define URAM288_BASE_ADDR_N  26
`define URAM288_BASE_ADDR_SZ 32
`define URAM288_BASE_DATA_SZ 144

// Attribute addresses
//

`define URAM288_BASE__AUTO_SLEEP_LATENCY    32'h00000000
`define URAM288_BASE__AUTO_SLEEP_LATENCY_SZ 32

`define URAM288_BASE__AVG_CONS_INACTIVE_CYCLES    32'h00000001
`define URAM288_BASE__AVG_CONS_INACTIVE_CYCLES_SZ 32

`define URAM288_BASE__BWE_MODE_A    32'h00000002
`define URAM288_BASE__BWE_MODE_A_SZ 144

`define URAM288_BASE__BWE_MODE_B    32'h00000003
`define URAM288_BASE__BWE_MODE_B_SZ 144

`define URAM288_BASE__EN_AUTO_SLEEP_MODE    32'h00000004
`define URAM288_BASE__EN_AUTO_SLEEP_MODE_SZ 40

`define URAM288_BASE__EN_ECC_RD_A    32'h00000005
`define URAM288_BASE__EN_ECC_RD_A_SZ 40

`define URAM288_BASE__EN_ECC_RD_B    32'h00000006
`define URAM288_BASE__EN_ECC_RD_B_SZ 40

`define URAM288_BASE__EN_ECC_WR_A    32'h00000007
`define URAM288_BASE__EN_ECC_WR_A_SZ 40

`define URAM288_BASE__EN_ECC_WR_B    32'h00000008
`define URAM288_BASE__EN_ECC_WR_B_SZ 40

`define URAM288_BASE__IREG_PRE_A    32'h00000009
`define URAM288_BASE__IREG_PRE_A_SZ 40

`define URAM288_BASE__IREG_PRE_B    32'h0000000a
`define URAM288_BASE__IREG_PRE_B_SZ 40

`define URAM288_BASE__IS_CLK_INVERTED    32'h0000000b
`define URAM288_BASE__IS_CLK_INVERTED_SZ 1

`define URAM288_BASE__IS_EN_A_INVERTED    32'h0000000c
`define URAM288_BASE__IS_EN_A_INVERTED_SZ 1

`define URAM288_BASE__IS_EN_B_INVERTED    32'h0000000d
`define URAM288_BASE__IS_EN_B_INVERTED_SZ 1

`define URAM288_BASE__IS_RDB_WR_A_INVERTED    32'h0000000e
`define URAM288_BASE__IS_RDB_WR_A_INVERTED_SZ 1

`define URAM288_BASE__IS_RDB_WR_B_INVERTED    32'h0000000f
`define URAM288_BASE__IS_RDB_WR_B_INVERTED_SZ 1

`define URAM288_BASE__IS_RST_A_INVERTED    32'h00000010
`define URAM288_BASE__IS_RST_A_INVERTED_SZ 1

`define URAM288_BASE__IS_RST_B_INVERTED    32'h00000011
`define URAM288_BASE__IS_RST_B_INVERTED_SZ 1

`define URAM288_BASE__OREG_A    32'h00000012
`define URAM288_BASE__OREG_A_SZ 40

`define URAM288_BASE__OREG_B    32'h00000013
`define URAM288_BASE__OREG_B_SZ 40

`define URAM288_BASE__OREG_ECC_A    32'h00000014
`define URAM288_BASE__OREG_ECC_A_SZ 40

`define URAM288_BASE__OREG_ECC_B    32'h00000015
`define URAM288_BASE__OREG_ECC_B_SZ 40

`define URAM288_BASE__RST_MODE_A    32'h00000016
`define URAM288_BASE__RST_MODE_A_SZ 40

`define URAM288_BASE__RST_MODE_B    32'h00000017
`define URAM288_BASE__RST_MODE_B_SZ 40

`define URAM288_BASE__USE_EXT_CE_A    32'h00000018
`define URAM288_BASE__USE_EXT_CE_A_SZ 40

`define URAM288_BASE__USE_EXT_CE_B    32'h00000019
`define URAM288_BASE__USE_EXT_CE_B_SZ 40

`endif  // B_URAM288_BASE_DEFINES_VH