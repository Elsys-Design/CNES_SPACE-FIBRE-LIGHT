// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_IOBUFDS_COMP_DEFINES_VH
`else
`define B_IOBUFDS_COMP_DEFINES_VH

// Look-up table parameters
//

`define IOBUFDS_COMP_ADDR_N  4
`define IOBUFDS_COMP_ADDR_SZ 32
`define IOBUFDS_COMP_DATA_SZ 72

// Attribute addresses
//

`define IOBUFDS_COMP__DQS_BIAS    32'h00000000
`define IOBUFDS_COMP__DQS_BIAS_SZ 40

`define IOBUFDS_COMP__IBUF_LOW_PWR    32'h00000001
`define IOBUFDS_COMP__IBUF_LOW_PWR_SZ 40

`define IOBUFDS_COMP__IOSTANDARD    32'h00000002
`define IOBUFDS_COMP__IOSTANDARD_SZ 56

`define IOBUFDS_COMP__USE_IBUFDISABLE    32'h00000003
`define IOBUFDS_COMP__USE_IBUFDISABLE_SZ 72

`endif  // B_IOBUFDS_COMP_DEFINES_VH