// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_HBM_TWO_STACK_INTF_DEFINES_VH
`else
`define B_HBM_TWO_STACK_INTF_DEFINES_VH

// Look-up table parameters
//

`define HBM_TWO_STACK_INTF_ADDR_N  241
`define HBM_TWO_STACK_INTF_ADDR_SZ 32
`define HBM_TWO_STACK_INTF_DATA_SZ 152

// Attribute addresses
//

`define HBM_TWO_STACK_INTF__CLK_SEL_00    32'h00000000
`define HBM_TWO_STACK_INTF__CLK_SEL_00_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_01    32'h00000001
`define HBM_TWO_STACK_INTF__CLK_SEL_01_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_02    32'h00000002
`define HBM_TWO_STACK_INTF__CLK_SEL_02_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_03    32'h00000003
`define HBM_TWO_STACK_INTF__CLK_SEL_03_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_04    32'h00000004
`define HBM_TWO_STACK_INTF__CLK_SEL_04_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_05    32'h00000005
`define HBM_TWO_STACK_INTF__CLK_SEL_05_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_06    32'h00000006
`define HBM_TWO_STACK_INTF__CLK_SEL_06_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_07    32'h00000007
`define HBM_TWO_STACK_INTF__CLK_SEL_07_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_08    32'h00000008
`define HBM_TWO_STACK_INTF__CLK_SEL_08_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_09    32'h00000009
`define HBM_TWO_STACK_INTF__CLK_SEL_09_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_10    32'h0000000a
`define HBM_TWO_STACK_INTF__CLK_SEL_10_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_11    32'h0000000b
`define HBM_TWO_STACK_INTF__CLK_SEL_11_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_12    32'h0000000c
`define HBM_TWO_STACK_INTF__CLK_SEL_12_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_13    32'h0000000d
`define HBM_TWO_STACK_INTF__CLK_SEL_13_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_14    32'h0000000e
`define HBM_TWO_STACK_INTF__CLK_SEL_14_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_15    32'h0000000f
`define HBM_TWO_STACK_INTF__CLK_SEL_15_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_16    32'h00000010
`define HBM_TWO_STACK_INTF__CLK_SEL_16_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_17    32'h00000011
`define HBM_TWO_STACK_INTF__CLK_SEL_17_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_18    32'h00000012
`define HBM_TWO_STACK_INTF__CLK_SEL_18_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_19    32'h00000013
`define HBM_TWO_STACK_INTF__CLK_SEL_19_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_20    32'h00000014
`define HBM_TWO_STACK_INTF__CLK_SEL_20_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_21    32'h00000015
`define HBM_TWO_STACK_INTF__CLK_SEL_21_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_22    32'h00000016
`define HBM_TWO_STACK_INTF__CLK_SEL_22_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_23    32'h00000017
`define HBM_TWO_STACK_INTF__CLK_SEL_23_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_24    32'h00000018
`define HBM_TWO_STACK_INTF__CLK_SEL_24_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_25    32'h00000019
`define HBM_TWO_STACK_INTF__CLK_SEL_25_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_26    32'h0000001a
`define HBM_TWO_STACK_INTF__CLK_SEL_26_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_27    32'h0000001b
`define HBM_TWO_STACK_INTF__CLK_SEL_27_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_28    32'h0000001c
`define HBM_TWO_STACK_INTF__CLK_SEL_28_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_29    32'h0000001d
`define HBM_TWO_STACK_INTF__CLK_SEL_29_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_30    32'h0000001e
`define HBM_TWO_STACK_INTF__CLK_SEL_30_SZ 40

`define HBM_TWO_STACK_INTF__CLK_SEL_31    32'h0000001f
`define HBM_TWO_STACK_INTF__CLK_SEL_31_SZ 40

`define HBM_TWO_STACK_INTF__DATARATE_00    32'h00000020
`define HBM_TWO_STACK_INTF__DATARATE_00_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_01    32'h00000021
`define HBM_TWO_STACK_INTF__DATARATE_01_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_02    32'h00000022
`define HBM_TWO_STACK_INTF__DATARATE_02_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_03    32'h00000023
`define HBM_TWO_STACK_INTF__DATARATE_03_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_04    32'h00000024
`define HBM_TWO_STACK_INTF__DATARATE_04_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_05    32'h00000025
`define HBM_TWO_STACK_INTF__DATARATE_05_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_06    32'h00000026
`define HBM_TWO_STACK_INTF__DATARATE_06_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_07    32'h00000027
`define HBM_TWO_STACK_INTF__DATARATE_07_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_08    32'h00000028
`define HBM_TWO_STACK_INTF__DATARATE_08_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_09    32'h00000029
`define HBM_TWO_STACK_INTF__DATARATE_09_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_10    32'h0000002a
`define HBM_TWO_STACK_INTF__DATARATE_10_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_11    32'h0000002b
`define HBM_TWO_STACK_INTF__DATARATE_11_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_12    32'h0000002c
`define HBM_TWO_STACK_INTF__DATARATE_12_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_13    32'h0000002d
`define HBM_TWO_STACK_INTF__DATARATE_13_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_14    32'h0000002e
`define HBM_TWO_STACK_INTF__DATARATE_14_SZ 11

`define HBM_TWO_STACK_INTF__DATARATE_15    32'h0000002f
`define HBM_TWO_STACK_INTF__DATARATE_15_SZ 11

`define HBM_TWO_STACK_INTF__DA_LOCKOUT_0    32'h00000030
`define HBM_TWO_STACK_INTF__DA_LOCKOUT_0_SZ 40

`define HBM_TWO_STACK_INTF__DA_LOCKOUT_1    32'h00000031
`define HBM_TWO_STACK_INTF__DA_LOCKOUT_1_SZ 40

`define HBM_TWO_STACK_INTF__IS_APB_0_PCLK_INVERTED    32'h00000032
`define HBM_TWO_STACK_INTF__IS_APB_0_PCLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_APB_0_PRESET_N_INVERTED    32'h00000033
`define HBM_TWO_STACK_INTF__IS_APB_0_PRESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_APB_1_PCLK_INVERTED    32'h00000034
`define HBM_TWO_STACK_INTF__IS_APB_1_PCLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_APB_1_PRESET_N_INVERTED    32'h00000035
`define HBM_TWO_STACK_INTF__IS_APB_1_PRESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_00_ACLK_INVERTED    32'h00000036
`define HBM_TWO_STACK_INTF__IS_AXI_00_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_00_ARESET_N_INVERTED    32'h00000037
`define HBM_TWO_STACK_INTF__IS_AXI_00_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_01_ACLK_INVERTED    32'h00000038
`define HBM_TWO_STACK_INTF__IS_AXI_01_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_01_ARESET_N_INVERTED    32'h00000039
`define HBM_TWO_STACK_INTF__IS_AXI_01_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_02_ACLK_INVERTED    32'h0000003a
`define HBM_TWO_STACK_INTF__IS_AXI_02_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_02_ARESET_N_INVERTED    32'h0000003b
`define HBM_TWO_STACK_INTF__IS_AXI_02_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_03_ACLK_INVERTED    32'h0000003c
`define HBM_TWO_STACK_INTF__IS_AXI_03_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_03_ARESET_N_INVERTED    32'h0000003d
`define HBM_TWO_STACK_INTF__IS_AXI_03_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_04_ACLK_INVERTED    32'h0000003e
`define HBM_TWO_STACK_INTF__IS_AXI_04_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_04_ARESET_N_INVERTED    32'h0000003f
`define HBM_TWO_STACK_INTF__IS_AXI_04_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_05_ACLK_INVERTED    32'h00000040
`define HBM_TWO_STACK_INTF__IS_AXI_05_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_05_ARESET_N_INVERTED    32'h00000041
`define HBM_TWO_STACK_INTF__IS_AXI_05_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_06_ACLK_INVERTED    32'h00000042
`define HBM_TWO_STACK_INTF__IS_AXI_06_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_06_ARESET_N_INVERTED    32'h00000043
`define HBM_TWO_STACK_INTF__IS_AXI_06_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_07_ACLK_INVERTED    32'h00000044
`define HBM_TWO_STACK_INTF__IS_AXI_07_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_07_ARESET_N_INVERTED    32'h00000045
`define HBM_TWO_STACK_INTF__IS_AXI_07_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_08_ACLK_INVERTED    32'h00000046
`define HBM_TWO_STACK_INTF__IS_AXI_08_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_08_ARESET_N_INVERTED    32'h00000047
`define HBM_TWO_STACK_INTF__IS_AXI_08_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_09_ACLK_INVERTED    32'h00000048
`define HBM_TWO_STACK_INTF__IS_AXI_09_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_09_ARESET_N_INVERTED    32'h00000049
`define HBM_TWO_STACK_INTF__IS_AXI_09_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_10_ACLK_INVERTED    32'h0000004a
`define HBM_TWO_STACK_INTF__IS_AXI_10_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_10_ARESET_N_INVERTED    32'h0000004b
`define HBM_TWO_STACK_INTF__IS_AXI_10_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_11_ACLK_INVERTED    32'h0000004c
`define HBM_TWO_STACK_INTF__IS_AXI_11_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_11_ARESET_N_INVERTED    32'h0000004d
`define HBM_TWO_STACK_INTF__IS_AXI_11_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_12_ACLK_INVERTED    32'h0000004e
`define HBM_TWO_STACK_INTF__IS_AXI_12_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_12_ARESET_N_INVERTED    32'h0000004f
`define HBM_TWO_STACK_INTF__IS_AXI_12_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_13_ACLK_INVERTED    32'h00000050
`define HBM_TWO_STACK_INTF__IS_AXI_13_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_13_ARESET_N_INVERTED    32'h00000051
`define HBM_TWO_STACK_INTF__IS_AXI_13_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_14_ACLK_INVERTED    32'h00000052
`define HBM_TWO_STACK_INTF__IS_AXI_14_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_14_ARESET_N_INVERTED    32'h00000053
`define HBM_TWO_STACK_INTF__IS_AXI_14_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_15_ACLK_INVERTED    32'h00000054
`define HBM_TWO_STACK_INTF__IS_AXI_15_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_15_ARESET_N_INVERTED    32'h00000055
`define HBM_TWO_STACK_INTF__IS_AXI_15_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_16_ACLK_INVERTED    32'h00000056
`define HBM_TWO_STACK_INTF__IS_AXI_16_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_16_ARESET_N_INVERTED    32'h00000057
`define HBM_TWO_STACK_INTF__IS_AXI_16_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_17_ACLK_INVERTED    32'h00000058
`define HBM_TWO_STACK_INTF__IS_AXI_17_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_17_ARESET_N_INVERTED    32'h00000059
`define HBM_TWO_STACK_INTF__IS_AXI_17_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_18_ACLK_INVERTED    32'h0000005a
`define HBM_TWO_STACK_INTF__IS_AXI_18_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_18_ARESET_N_INVERTED    32'h0000005b
`define HBM_TWO_STACK_INTF__IS_AXI_18_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_19_ACLK_INVERTED    32'h0000005c
`define HBM_TWO_STACK_INTF__IS_AXI_19_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_19_ARESET_N_INVERTED    32'h0000005d
`define HBM_TWO_STACK_INTF__IS_AXI_19_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_20_ACLK_INVERTED    32'h0000005e
`define HBM_TWO_STACK_INTF__IS_AXI_20_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_20_ARESET_N_INVERTED    32'h0000005f
`define HBM_TWO_STACK_INTF__IS_AXI_20_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_21_ACLK_INVERTED    32'h00000060
`define HBM_TWO_STACK_INTF__IS_AXI_21_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_21_ARESET_N_INVERTED    32'h00000061
`define HBM_TWO_STACK_INTF__IS_AXI_21_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_22_ACLK_INVERTED    32'h00000062
`define HBM_TWO_STACK_INTF__IS_AXI_22_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_22_ARESET_N_INVERTED    32'h00000063
`define HBM_TWO_STACK_INTF__IS_AXI_22_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_23_ACLK_INVERTED    32'h00000064
`define HBM_TWO_STACK_INTF__IS_AXI_23_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_23_ARESET_N_INVERTED    32'h00000065
`define HBM_TWO_STACK_INTF__IS_AXI_23_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_24_ACLK_INVERTED    32'h00000066
`define HBM_TWO_STACK_INTF__IS_AXI_24_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_24_ARESET_N_INVERTED    32'h00000067
`define HBM_TWO_STACK_INTF__IS_AXI_24_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_25_ACLK_INVERTED    32'h00000068
`define HBM_TWO_STACK_INTF__IS_AXI_25_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_25_ARESET_N_INVERTED    32'h00000069
`define HBM_TWO_STACK_INTF__IS_AXI_25_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_26_ACLK_INVERTED    32'h0000006a
`define HBM_TWO_STACK_INTF__IS_AXI_26_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_26_ARESET_N_INVERTED    32'h0000006b
`define HBM_TWO_STACK_INTF__IS_AXI_26_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_27_ACLK_INVERTED    32'h0000006c
`define HBM_TWO_STACK_INTF__IS_AXI_27_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_27_ARESET_N_INVERTED    32'h0000006d
`define HBM_TWO_STACK_INTF__IS_AXI_27_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_28_ACLK_INVERTED    32'h0000006e
`define HBM_TWO_STACK_INTF__IS_AXI_28_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_28_ARESET_N_INVERTED    32'h0000006f
`define HBM_TWO_STACK_INTF__IS_AXI_28_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_29_ACLK_INVERTED    32'h00000070
`define HBM_TWO_STACK_INTF__IS_AXI_29_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_29_ARESET_N_INVERTED    32'h00000071
`define HBM_TWO_STACK_INTF__IS_AXI_29_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_30_ACLK_INVERTED    32'h00000072
`define HBM_TWO_STACK_INTF__IS_AXI_30_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_30_ARESET_N_INVERTED    32'h00000073
`define HBM_TWO_STACK_INTF__IS_AXI_30_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_31_ACLK_INVERTED    32'h00000074
`define HBM_TWO_STACK_INTF__IS_AXI_31_ACLK_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__IS_AXI_31_ARESET_N_INVERTED    32'h00000075
`define HBM_TWO_STACK_INTF__IS_AXI_31_ARESET_N_INVERTED_SZ 1

`define HBM_TWO_STACK_INTF__MC_ENABLE_00    32'h00000076
`define HBM_TWO_STACK_INTF__MC_ENABLE_00_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_01    32'h00000077
`define HBM_TWO_STACK_INTF__MC_ENABLE_01_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_02    32'h00000078
`define HBM_TWO_STACK_INTF__MC_ENABLE_02_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_03    32'h00000079
`define HBM_TWO_STACK_INTF__MC_ENABLE_03_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_04    32'h0000007a
`define HBM_TWO_STACK_INTF__MC_ENABLE_04_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_05    32'h0000007b
`define HBM_TWO_STACK_INTF__MC_ENABLE_05_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_06    32'h0000007c
`define HBM_TWO_STACK_INTF__MC_ENABLE_06_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_07    32'h0000007d
`define HBM_TWO_STACK_INTF__MC_ENABLE_07_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_08    32'h0000007e
`define HBM_TWO_STACK_INTF__MC_ENABLE_08_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_09    32'h0000007f
`define HBM_TWO_STACK_INTF__MC_ENABLE_09_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_10    32'h00000080
`define HBM_TWO_STACK_INTF__MC_ENABLE_10_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_11    32'h00000081
`define HBM_TWO_STACK_INTF__MC_ENABLE_11_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_12    32'h00000082
`define HBM_TWO_STACK_INTF__MC_ENABLE_12_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_13    32'h00000083
`define HBM_TWO_STACK_INTF__MC_ENABLE_13_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_14    32'h00000084
`define HBM_TWO_STACK_INTF__MC_ENABLE_14_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_15    32'h00000085
`define HBM_TWO_STACK_INTF__MC_ENABLE_15_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_APB_00    32'h00000086
`define HBM_TWO_STACK_INTF__MC_ENABLE_APB_00_SZ 40

`define HBM_TWO_STACK_INTF__MC_ENABLE_APB_01    32'h00000087
`define HBM_TWO_STACK_INTF__MC_ENABLE_APB_01_SZ 40

`define HBM_TWO_STACK_INTF__PAGEHIT_PERCENT_00    32'h00000088
`define HBM_TWO_STACK_INTF__PAGEHIT_PERCENT_00_SZ 7

`define HBM_TWO_STACK_INTF__PAGEHIT_PERCENT_01    32'h00000089
`define HBM_TWO_STACK_INTF__PAGEHIT_PERCENT_01_SZ 7

`define HBM_TWO_STACK_INTF__PHY_ENABLE_00    32'h0000008a
`define HBM_TWO_STACK_INTF__PHY_ENABLE_00_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_01    32'h0000008b
`define HBM_TWO_STACK_INTF__PHY_ENABLE_01_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_02    32'h0000008c
`define HBM_TWO_STACK_INTF__PHY_ENABLE_02_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_03    32'h0000008d
`define HBM_TWO_STACK_INTF__PHY_ENABLE_03_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_04    32'h0000008e
`define HBM_TWO_STACK_INTF__PHY_ENABLE_04_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_05    32'h0000008f
`define HBM_TWO_STACK_INTF__PHY_ENABLE_05_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_06    32'h00000090
`define HBM_TWO_STACK_INTF__PHY_ENABLE_06_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_07    32'h00000091
`define HBM_TWO_STACK_INTF__PHY_ENABLE_07_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_08    32'h00000092
`define HBM_TWO_STACK_INTF__PHY_ENABLE_08_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_09    32'h00000093
`define HBM_TWO_STACK_INTF__PHY_ENABLE_09_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_10    32'h00000094
`define HBM_TWO_STACK_INTF__PHY_ENABLE_10_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_11    32'h00000095
`define HBM_TWO_STACK_INTF__PHY_ENABLE_11_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_12    32'h00000096
`define HBM_TWO_STACK_INTF__PHY_ENABLE_12_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_13    32'h00000097
`define HBM_TWO_STACK_INTF__PHY_ENABLE_13_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_14    32'h00000098
`define HBM_TWO_STACK_INTF__PHY_ENABLE_14_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_15    32'h00000099
`define HBM_TWO_STACK_INTF__PHY_ENABLE_15_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_16    32'h0000009a
`define HBM_TWO_STACK_INTF__PHY_ENABLE_16_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_17    32'h0000009b
`define HBM_TWO_STACK_INTF__PHY_ENABLE_17_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_18    32'h0000009c
`define HBM_TWO_STACK_INTF__PHY_ENABLE_18_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_19    32'h0000009d
`define HBM_TWO_STACK_INTF__PHY_ENABLE_19_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_20    32'h0000009e
`define HBM_TWO_STACK_INTF__PHY_ENABLE_20_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_21    32'h0000009f
`define HBM_TWO_STACK_INTF__PHY_ENABLE_21_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_22    32'h000000a0
`define HBM_TWO_STACK_INTF__PHY_ENABLE_22_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_23    32'h000000a1
`define HBM_TWO_STACK_INTF__PHY_ENABLE_23_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_24    32'h000000a2
`define HBM_TWO_STACK_INTF__PHY_ENABLE_24_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_25    32'h000000a3
`define HBM_TWO_STACK_INTF__PHY_ENABLE_25_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_26    32'h000000a4
`define HBM_TWO_STACK_INTF__PHY_ENABLE_26_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_27    32'h000000a5
`define HBM_TWO_STACK_INTF__PHY_ENABLE_27_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_28    32'h000000a6
`define HBM_TWO_STACK_INTF__PHY_ENABLE_28_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_29    32'h000000a7
`define HBM_TWO_STACK_INTF__PHY_ENABLE_29_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_30    32'h000000a8
`define HBM_TWO_STACK_INTF__PHY_ENABLE_30_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_31    32'h000000a9
`define HBM_TWO_STACK_INTF__PHY_ENABLE_31_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_APB_00    32'h000000aa
`define HBM_TWO_STACK_INTF__PHY_ENABLE_APB_00_SZ 40

`define HBM_TWO_STACK_INTF__PHY_ENABLE_APB_01    32'h000000ab
`define HBM_TWO_STACK_INTF__PHY_ENABLE_APB_01_SZ 40

`define HBM_TWO_STACK_INTF__PHY_PCLK_INVERT_01    32'h000000ac
`define HBM_TWO_STACK_INTF__PHY_PCLK_INVERT_01_SZ 40

`define HBM_TWO_STACK_INTF__PHY_PCLK_INVERT_02    32'h000000ad
`define HBM_TWO_STACK_INTF__PHY_PCLK_INVERT_02_SZ 40

`define HBM_TWO_STACK_INTF__READ_PERCENT_00    32'h000000ae
`define HBM_TWO_STACK_INTF__READ_PERCENT_00_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_01    32'h000000af
`define HBM_TWO_STACK_INTF__READ_PERCENT_01_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_02    32'h000000b0
`define HBM_TWO_STACK_INTF__READ_PERCENT_02_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_03    32'h000000b1
`define HBM_TWO_STACK_INTF__READ_PERCENT_03_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_04    32'h000000b2
`define HBM_TWO_STACK_INTF__READ_PERCENT_04_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_05    32'h000000b3
`define HBM_TWO_STACK_INTF__READ_PERCENT_05_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_06    32'h000000b4
`define HBM_TWO_STACK_INTF__READ_PERCENT_06_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_07    32'h000000b5
`define HBM_TWO_STACK_INTF__READ_PERCENT_07_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_08    32'h000000b6
`define HBM_TWO_STACK_INTF__READ_PERCENT_08_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_09    32'h000000b7
`define HBM_TWO_STACK_INTF__READ_PERCENT_09_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_10    32'h000000b8
`define HBM_TWO_STACK_INTF__READ_PERCENT_10_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_11    32'h000000b9
`define HBM_TWO_STACK_INTF__READ_PERCENT_11_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_12    32'h000000ba
`define HBM_TWO_STACK_INTF__READ_PERCENT_12_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_13    32'h000000bb
`define HBM_TWO_STACK_INTF__READ_PERCENT_13_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_14    32'h000000bc
`define HBM_TWO_STACK_INTF__READ_PERCENT_14_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_15    32'h000000bd
`define HBM_TWO_STACK_INTF__READ_PERCENT_15_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_16    32'h000000be
`define HBM_TWO_STACK_INTF__READ_PERCENT_16_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_17    32'h000000bf
`define HBM_TWO_STACK_INTF__READ_PERCENT_17_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_18    32'h000000c0
`define HBM_TWO_STACK_INTF__READ_PERCENT_18_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_19    32'h000000c1
`define HBM_TWO_STACK_INTF__READ_PERCENT_19_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_20    32'h000000c2
`define HBM_TWO_STACK_INTF__READ_PERCENT_20_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_21    32'h000000c3
`define HBM_TWO_STACK_INTF__READ_PERCENT_21_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_22    32'h000000c4
`define HBM_TWO_STACK_INTF__READ_PERCENT_22_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_23    32'h000000c5
`define HBM_TWO_STACK_INTF__READ_PERCENT_23_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_24    32'h000000c6
`define HBM_TWO_STACK_INTF__READ_PERCENT_24_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_25    32'h000000c7
`define HBM_TWO_STACK_INTF__READ_PERCENT_25_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_26    32'h000000c8
`define HBM_TWO_STACK_INTF__READ_PERCENT_26_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_27    32'h000000c9
`define HBM_TWO_STACK_INTF__READ_PERCENT_27_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_28    32'h000000ca
`define HBM_TWO_STACK_INTF__READ_PERCENT_28_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_29    32'h000000cb
`define HBM_TWO_STACK_INTF__READ_PERCENT_29_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_30    32'h000000cc
`define HBM_TWO_STACK_INTF__READ_PERCENT_30_SZ 7

`define HBM_TWO_STACK_INTF__READ_PERCENT_31    32'h000000cd
`define HBM_TWO_STACK_INTF__READ_PERCENT_31_SZ 7

`define HBM_TWO_STACK_INTF__SIM_DEVICE    32'h000000ce
`define HBM_TWO_STACK_INTF__SIM_DEVICE_SZ 152

`define HBM_TWO_STACK_INTF__SWITCH_ENABLE_00    32'h000000cf
`define HBM_TWO_STACK_INTF__SWITCH_ENABLE_00_SZ 40

`define HBM_TWO_STACK_INTF__SWITCH_ENABLE_01    32'h000000d0
`define HBM_TWO_STACK_INTF__SWITCH_ENABLE_01_SZ 40

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_00    32'h000000d1
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_00_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_01    32'h000000d2
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_01_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_02    32'h000000d3
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_02_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_03    32'h000000d4
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_03_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_04    32'h000000d5
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_04_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_05    32'h000000d6
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_05_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_06    32'h000000d7
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_06_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_07    32'h000000d8
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_07_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_08    32'h000000d9
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_08_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_09    32'h000000da
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_09_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_10    32'h000000db
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_10_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_11    32'h000000dc
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_11_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_12    32'h000000dd
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_12_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_13    32'h000000de
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_13_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_14    32'h000000df
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_14_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_15    32'h000000e0
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_15_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_16    32'h000000e1
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_16_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_17    32'h000000e2
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_17_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_18    32'h000000e3
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_18_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_19    32'h000000e4
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_19_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_20    32'h000000e5
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_20_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_21    32'h000000e6
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_21_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_22    32'h000000e7
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_22_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_23    32'h000000e8
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_23_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_24    32'h000000e9
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_24_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_25    32'h000000ea
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_25_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_26    32'h000000eb
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_26_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_27    32'h000000ec
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_27_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_28    32'h000000ed
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_28_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_29    32'h000000ee
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_29_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_30    32'h000000ef
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_30_SZ 7

`define HBM_TWO_STACK_INTF__WRITE_PERCENT_31    32'h000000f0
`define HBM_TWO_STACK_INTF__WRITE_PERCENT_31_SZ 7

`endif  // B_HBM_TWO_STACK_INTF_DEFINES_VH