// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_MBUFGCTRL_DEFINES_VH
`else
`define B_MBUFGCTRL_DEFINES_VH

// Look-up table parameters
//

`define MBUFGCTRL_ADDR_N  16
`define MBUFGCTRL_ADDR_SZ 32
`define MBUFGCTRL_DATA_SZ 144

// Attribute addresses
//

`define MBUFGCTRL__CE_TYPE_CE0    32'h00000000
`define MBUFGCTRL__CE_TYPE_CE0_SZ 64

`define MBUFGCTRL__CE_TYPE_CE1    32'h00000001
`define MBUFGCTRL__CE_TYPE_CE1_SZ 64

`define MBUFGCTRL__INIT_OUT    32'h00000002
`define MBUFGCTRL__INIT_OUT_SZ 32

`define MBUFGCTRL__IS_CE0_INVERTED    32'h00000003
`define MBUFGCTRL__IS_CE0_INVERTED_SZ 1

`define MBUFGCTRL__IS_CE1_INVERTED    32'h00000004
`define MBUFGCTRL__IS_CE1_INVERTED_SZ 1

`define MBUFGCTRL__IS_I0_INVERTED    32'h00000005
`define MBUFGCTRL__IS_I0_INVERTED_SZ 1

`define MBUFGCTRL__IS_I1_INVERTED    32'h00000006
`define MBUFGCTRL__IS_I1_INVERTED_SZ 1

`define MBUFGCTRL__IS_IGNORE0_INVERTED    32'h00000007
`define MBUFGCTRL__IS_IGNORE0_INVERTED_SZ 1

`define MBUFGCTRL__IS_IGNORE1_INVERTED    32'h00000008
`define MBUFGCTRL__IS_IGNORE1_INVERTED_SZ 1

`define MBUFGCTRL__IS_S0_INVERTED    32'h00000009
`define MBUFGCTRL__IS_S0_INVERTED_SZ 1

`define MBUFGCTRL__IS_S1_INVERTED    32'h0000000a
`define MBUFGCTRL__IS_S1_INVERTED_SZ 1

`define MBUFGCTRL__MODE    32'h0000000b
`define MBUFGCTRL__MODE_SZ 88

`define MBUFGCTRL__PRESELECT_I0    32'h0000000c
`define MBUFGCTRL__PRESELECT_I0_SZ 40

`define MBUFGCTRL__PRESELECT_I1    32'h0000000d
`define MBUFGCTRL__PRESELECT_I1_SZ 40

`define MBUFGCTRL__SIM_DEVICE    32'h0000000e
`define MBUFGCTRL__SIM_DEVICE_SZ 144

`define MBUFGCTRL__STARTUP_SYNC    32'h0000000f
`define MBUFGCTRL__STARTUP_SYNC_SZ 40

`endif  // B_MBUFGCTRL_DEFINES_VH
