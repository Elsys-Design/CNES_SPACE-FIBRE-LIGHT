// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_NOC2_NPS7575_DEFINES_VH
`else
`define B_NOC2_NPS7575_DEFINES_VH

// Look-up table parameters
//

`define NOC2_NPS7575_ADDR_N  195
`define NOC2_NPS7575_ADDR_SZ 32
`define NOC2_NPS7575_DATA_SZ 32

// Attribute addresses
//

`define NOC2_NPS7575__REG_CLOCK_MUX    32'h00000000
`define NOC2_NPS7575__REG_CLOCK_MUX_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID0_P01    32'h00000001
`define NOC2_NPS7575__REG_HIGH_ID0_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID0_P23    32'h00000002
`define NOC2_NPS7575__REG_HIGH_ID0_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID10_P01    32'h00000003
`define NOC2_NPS7575__REG_HIGH_ID10_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID10_P23    32'h00000004
`define NOC2_NPS7575__REG_HIGH_ID10_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID11_P01    32'h00000005
`define NOC2_NPS7575__REG_HIGH_ID11_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID11_P23    32'h00000006
`define NOC2_NPS7575__REG_HIGH_ID11_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID12_P01    32'h00000007
`define NOC2_NPS7575__REG_HIGH_ID12_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID12_P23    32'h00000008
`define NOC2_NPS7575__REG_HIGH_ID12_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID13_P01    32'h00000009
`define NOC2_NPS7575__REG_HIGH_ID13_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID13_P23    32'h0000000a
`define NOC2_NPS7575__REG_HIGH_ID13_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID14_P01    32'h0000000b
`define NOC2_NPS7575__REG_HIGH_ID14_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID14_P23    32'h0000000c
`define NOC2_NPS7575__REG_HIGH_ID14_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID15_P01    32'h0000000d
`define NOC2_NPS7575__REG_HIGH_ID15_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID15_P23    32'h0000000e
`define NOC2_NPS7575__REG_HIGH_ID15_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID16_P01    32'h0000000f
`define NOC2_NPS7575__REG_HIGH_ID16_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID16_P23    32'h00000010
`define NOC2_NPS7575__REG_HIGH_ID16_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID17_P01    32'h00000011
`define NOC2_NPS7575__REG_HIGH_ID17_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID17_P23    32'h00000012
`define NOC2_NPS7575__REG_HIGH_ID17_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID18_P01    32'h00000013
`define NOC2_NPS7575__REG_HIGH_ID18_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID18_P23    32'h00000014
`define NOC2_NPS7575__REG_HIGH_ID18_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID19_P01    32'h00000015
`define NOC2_NPS7575__REG_HIGH_ID19_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID19_P23    32'h00000016
`define NOC2_NPS7575__REG_HIGH_ID19_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID1_P01    32'h00000017
`define NOC2_NPS7575__REG_HIGH_ID1_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID1_P23    32'h00000018
`define NOC2_NPS7575__REG_HIGH_ID1_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID20_P01    32'h00000019
`define NOC2_NPS7575__REG_HIGH_ID20_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID20_P23    32'h0000001a
`define NOC2_NPS7575__REG_HIGH_ID20_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID21_P01    32'h0000001b
`define NOC2_NPS7575__REG_HIGH_ID21_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID21_P23    32'h0000001c
`define NOC2_NPS7575__REG_HIGH_ID21_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID22_P01    32'h0000001d
`define NOC2_NPS7575__REG_HIGH_ID22_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID22_P23    32'h0000001e
`define NOC2_NPS7575__REG_HIGH_ID22_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID23_P01    32'h0000001f
`define NOC2_NPS7575__REG_HIGH_ID23_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID23_P23    32'h00000020
`define NOC2_NPS7575__REG_HIGH_ID23_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID24_P01    32'h00000021
`define NOC2_NPS7575__REG_HIGH_ID24_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID24_P23    32'h00000022
`define NOC2_NPS7575__REG_HIGH_ID24_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID25_P01    32'h00000023
`define NOC2_NPS7575__REG_HIGH_ID25_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID25_P23    32'h00000024
`define NOC2_NPS7575__REG_HIGH_ID25_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID26_P01    32'h00000025
`define NOC2_NPS7575__REG_HIGH_ID26_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID26_P23    32'h00000026
`define NOC2_NPS7575__REG_HIGH_ID26_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID27_P01    32'h00000027
`define NOC2_NPS7575__REG_HIGH_ID27_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID27_P23    32'h00000028
`define NOC2_NPS7575__REG_HIGH_ID27_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID28_P01    32'h00000029
`define NOC2_NPS7575__REG_HIGH_ID28_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID28_P23    32'h0000002a
`define NOC2_NPS7575__REG_HIGH_ID28_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID29_P01    32'h0000002b
`define NOC2_NPS7575__REG_HIGH_ID29_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID29_P23    32'h0000002c
`define NOC2_NPS7575__REG_HIGH_ID29_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID2_P01    32'h0000002d
`define NOC2_NPS7575__REG_HIGH_ID2_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID2_P23    32'h0000002e
`define NOC2_NPS7575__REG_HIGH_ID2_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID30_P01    32'h0000002f
`define NOC2_NPS7575__REG_HIGH_ID30_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID30_P23    32'h00000030
`define NOC2_NPS7575__REG_HIGH_ID30_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID31_P01    32'h00000031
`define NOC2_NPS7575__REG_HIGH_ID31_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID31_P23    32'h00000032
`define NOC2_NPS7575__REG_HIGH_ID31_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID32_P01    32'h00000033
`define NOC2_NPS7575__REG_HIGH_ID32_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID32_P23    32'h00000034
`define NOC2_NPS7575__REG_HIGH_ID32_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID33_P01    32'h00000035
`define NOC2_NPS7575__REG_HIGH_ID33_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID33_P23    32'h00000036
`define NOC2_NPS7575__REG_HIGH_ID33_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID34_P01    32'h00000037
`define NOC2_NPS7575__REG_HIGH_ID34_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID34_P23    32'h00000038
`define NOC2_NPS7575__REG_HIGH_ID34_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID35_P01    32'h00000039
`define NOC2_NPS7575__REG_HIGH_ID35_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID35_P23    32'h0000003a
`define NOC2_NPS7575__REG_HIGH_ID35_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID36_P01    32'h0000003b
`define NOC2_NPS7575__REG_HIGH_ID36_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID36_P23    32'h0000003c
`define NOC2_NPS7575__REG_HIGH_ID36_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID37_P01    32'h0000003d
`define NOC2_NPS7575__REG_HIGH_ID37_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID37_P23    32'h0000003e
`define NOC2_NPS7575__REG_HIGH_ID37_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID38_P01    32'h0000003f
`define NOC2_NPS7575__REG_HIGH_ID38_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID38_P23    32'h00000040
`define NOC2_NPS7575__REG_HIGH_ID38_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID39_P01    32'h00000041
`define NOC2_NPS7575__REG_HIGH_ID39_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID39_P23    32'h00000042
`define NOC2_NPS7575__REG_HIGH_ID39_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID3_P01    32'h00000043
`define NOC2_NPS7575__REG_HIGH_ID3_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID3_P23    32'h00000044
`define NOC2_NPS7575__REG_HIGH_ID3_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID40_P01    32'h00000045
`define NOC2_NPS7575__REG_HIGH_ID40_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID40_P23    32'h00000046
`define NOC2_NPS7575__REG_HIGH_ID40_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID41_P01    32'h00000047
`define NOC2_NPS7575__REG_HIGH_ID41_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID41_P23    32'h00000048
`define NOC2_NPS7575__REG_HIGH_ID41_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID42_P01    32'h00000049
`define NOC2_NPS7575__REG_HIGH_ID42_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID42_P23    32'h0000004a
`define NOC2_NPS7575__REG_HIGH_ID42_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID43_P01    32'h0000004b
`define NOC2_NPS7575__REG_HIGH_ID43_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID43_P23    32'h0000004c
`define NOC2_NPS7575__REG_HIGH_ID43_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID44_P01    32'h0000004d
`define NOC2_NPS7575__REG_HIGH_ID44_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID44_P23    32'h0000004e
`define NOC2_NPS7575__REG_HIGH_ID44_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID45_P01    32'h0000004f
`define NOC2_NPS7575__REG_HIGH_ID45_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID45_P23    32'h00000050
`define NOC2_NPS7575__REG_HIGH_ID45_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID46_P01    32'h00000051
`define NOC2_NPS7575__REG_HIGH_ID46_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID46_P23    32'h00000052
`define NOC2_NPS7575__REG_HIGH_ID46_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID47_P01    32'h00000053
`define NOC2_NPS7575__REG_HIGH_ID47_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID47_P23    32'h00000054
`define NOC2_NPS7575__REG_HIGH_ID47_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID48_P01    32'h00000055
`define NOC2_NPS7575__REG_HIGH_ID48_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID48_P23    32'h00000056
`define NOC2_NPS7575__REG_HIGH_ID48_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID49_P01    32'h00000057
`define NOC2_NPS7575__REG_HIGH_ID49_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID49_P23    32'h00000058
`define NOC2_NPS7575__REG_HIGH_ID49_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID4_P01    32'h00000059
`define NOC2_NPS7575__REG_HIGH_ID4_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID4_P23    32'h0000005a
`define NOC2_NPS7575__REG_HIGH_ID4_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID50_P01    32'h0000005b
`define NOC2_NPS7575__REG_HIGH_ID50_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID50_P23    32'h0000005c
`define NOC2_NPS7575__REG_HIGH_ID50_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID51_P01    32'h0000005d
`define NOC2_NPS7575__REG_HIGH_ID51_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID51_P23    32'h0000005e
`define NOC2_NPS7575__REG_HIGH_ID51_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID52_P01    32'h0000005f
`define NOC2_NPS7575__REG_HIGH_ID52_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID52_P23    32'h00000060
`define NOC2_NPS7575__REG_HIGH_ID52_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID53_P01    32'h00000061
`define NOC2_NPS7575__REG_HIGH_ID53_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID53_P23    32'h00000062
`define NOC2_NPS7575__REG_HIGH_ID53_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID54_P01    32'h00000063
`define NOC2_NPS7575__REG_HIGH_ID54_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID54_P23    32'h00000064
`define NOC2_NPS7575__REG_HIGH_ID54_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID55_P01    32'h00000065
`define NOC2_NPS7575__REG_HIGH_ID55_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID55_P23    32'h00000066
`define NOC2_NPS7575__REG_HIGH_ID55_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID56_P01    32'h00000067
`define NOC2_NPS7575__REG_HIGH_ID56_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID56_P23    32'h00000068
`define NOC2_NPS7575__REG_HIGH_ID56_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID57_P01    32'h00000069
`define NOC2_NPS7575__REG_HIGH_ID57_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID57_P23    32'h0000006a
`define NOC2_NPS7575__REG_HIGH_ID57_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID58_P01    32'h0000006b
`define NOC2_NPS7575__REG_HIGH_ID58_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID58_P23    32'h0000006c
`define NOC2_NPS7575__REG_HIGH_ID58_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID59_P01    32'h0000006d
`define NOC2_NPS7575__REG_HIGH_ID59_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID59_P23    32'h0000006e
`define NOC2_NPS7575__REG_HIGH_ID59_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID5_P01    32'h0000006f
`define NOC2_NPS7575__REG_HIGH_ID5_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID5_P23    32'h00000070
`define NOC2_NPS7575__REG_HIGH_ID5_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID60_P01    32'h00000071
`define NOC2_NPS7575__REG_HIGH_ID60_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID60_P23    32'h00000072
`define NOC2_NPS7575__REG_HIGH_ID60_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID61_P01    32'h00000073
`define NOC2_NPS7575__REG_HIGH_ID61_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID61_P23    32'h00000074
`define NOC2_NPS7575__REG_HIGH_ID61_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID62_P01    32'h00000075
`define NOC2_NPS7575__REG_HIGH_ID62_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID62_P23    32'h00000076
`define NOC2_NPS7575__REG_HIGH_ID62_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID63_P01    32'h00000077
`define NOC2_NPS7575__REG_HIGH_ID63_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID63_P23    32'h00000078
`define NOC2_NPS7575__REG_HIGH_ID63_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID6_P01    32'h00000079
`define NOC2_NPS7575__REG_HIGH_ID6_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID6_P23    32'h0000007a
`define NOC2_NPS7575__REG_HIGH_ID6_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID7_P01    32'h0000007b
`define NOC2_NPS7575__REG_HIGH_ID7_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID7_P23    32'h0000007c
`define NOC2_NPS7575__REG_HIGH_ID7_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID8_P01    32'h0000007d
`define NOC2_NPS7575__REG_HIGH_ID8_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID8_P23    32'h0000007e
`define NOC2_NPS7575__REG_HIGH_ID8_P23_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID9_P01    32'h0000007f
`define NOC2_NPS7575__REG_HIGH_ID9_P01_SZ 32

`define NOC2_NPS7575__REG_HIGH_ID9_P23    32'h00000080
`define NOC2_NPS7575__REG_HIGH_ID9_P23_SZ 32

`define NOC2_NPS7575__REG_ID    32'h00000081
`define NOC2_NPS7575__REG_ID_SZ 10

`define NOC2_NPS7575__REG_LOW_ID0_P01    32'h00000082
`define NOC2_NPS7575__REG_LOW_ID0_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID0_P23    32'h00000083
`define NOC2_NPS7575__REG_LOW_ID0_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID10_P01    32'h00000084
`define NOC2_NPS7575__REG_LOW_ID10_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID10_P23    32'h00000085
`define NOC2_NPS7575__REG_LOW_ID10_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID11_P01    32'h00000086
`define NOC2_NPS7575__REG_LOW_ID11_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID11_P23    32'h00000087
`define NOC2_NPS7575__REG_LOW_ID11_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID12_P01    32'h00000088
`define NOC2_NPS7575__REG_LOW_ID12_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID12_P23    32'h00000089
`define NOC2_NPS7575__REG_LOW_ID12_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID13_P01    32'h0000008a
`define NOC2_NPS7575__REG_LOW_ID13_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID13_P23    32'h0000008b
`define NOC2_NPS7575__REG_LOW_ID13_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID14_P01    32'h0000008c
`define NOC2_NPS7575__REG_LOW_ID14_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID14_P23    32'h0000008d
`define NOC2_NPS7575__REG_LOW_ID14_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID15_P01    32'h0000008e
`define NOC2_NPS7575__REG_LOW_ID15_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID15_P23    32'h0000008f
`define NOC2_NPS7575__REG_LOW_ID15_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID1_P01    32'h00000090
`define NOC2_NPS7575__REG_LOW_ID1_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID1_P23    32'h00000091
`define NOC2_NPS7575__REG_LOW_ID1_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID2_P01    32'h00000092
`define NOC2_NPS7575__REG_LOW_ID2_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID2_P23    32'h00000093
`define NOC2_NPS7575__REG_LOW_ID2_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID3_P01    32'h00000094
`define NOC2_NPS7575__REG_LOW_ID3_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID3_P23    32'h00000095
`define NOC2_NPS7575__REG_LOW_ID3_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID4_P01    32'h00000096
`define NOC2_NPS7575__REG_LOW_ID4_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID4_P23    32'h00000097
`define NOC2_NPS7575__REG_LOW_ID4_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID5_P01    32'h00000098
`define NOC2_NPS7575__REG_LOW_ID5_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID5_P23    32'h00000099
`define NOC2_NPS7575__REG_LOW_ID5_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID6_P01    32'h0000009a
`define NOC2_NPS7575__REG_LOW_ID6_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID6_P23    32'h0000009b
`define NOC2_NPS7575__REG_LOW_ID6_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID7_P01    32'h0000009c
`define NOC2_NPS7575__REG_LOW_ID7_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID7_P23    32'h0000009d
`define NOC2_NPS7575__REG_LOW_ID7_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID8_P01    32'h0000009e
`define NOC2_NPS7575__REG_LOW_ID8_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID8_P23    32'h0000009f
`define NOC2_NPS7575__REG_LOW_ID8_P23_SZ 32

`define NOC2_NPS7575__REG_LOW_ID9_P01    32'h000000a0
`define NOC2_NPS7575__REG_LOW_ID9_P01_SZ 32

`define NOC2_NPS7575__REG_LOW_ID9_P23    32'h000000a1
`define NOC2_NPS7575__REG_LOW_ID9_P23_SZ 32

`define NOC2_NPS7575__REG_MID_ID0_P01    32'h000000a2
`define NOC2_NPS7575__REG_MID_ID0_P01_SZ 32

`define NOC2_NPS7575__REG_MID_ID0_P23    32'h000000a3
`define NOC2_NPS7575__REG_MID_ID0_P23_SZ 32

`define NOC2_NPS7575__REG_MID_ID1_P01    32'h000000a4
`define NOC2_NPS7575__REG_MID_ID1_P01_SZ 32

`define NOC2_NPS7575__REG_MID_ID1_P23    32'h000000a5
`define NOC2_NPS7575__REG_MID_ID1_P23_SZ 32

`define NOC2_NPS7575__REG_MID_ID2_P01    32'h000000a6
`define NOC2_NPS7575__REG_MID_ID2_P01_SZ 32

`define NOC2_NPS7575__REG_MID_ID2_P23    32'h000000a7
`define NOC2_NPS7575__REG_MID_ID2_P23_SZ 32

`define NOC2_NPS7575__REG_MID_ID3_P01    32'h000000a8
`define NOC2_NPS7575__REG_MID_ID3_P01_SZ 32

`define NOC2_NPS7575__REG_MID_ID3_P23    32'h000000a9
`define NOC2_NPS7575__REG_MID_ID3_P23_SZ 32

`define NOC2_NPS7575__REG_NOC_CTL    32'h000000aa
`define NOC2_NPS7575__REG_NOC_CTL_SZ 16

`define NOC2_NPS7575__REG_P00_P1_0_VCA_TOKEN    32'h000000ab
`define NOC2_NPS7575__REG_P00_P1_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P00_P1_1_VCA_TOKEN    32'h000000ac
`define NOC2_NPS7575__REG_P00_P1_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P01_P2_0_VCA_TOKEN    32'h000000ad
`define NOC2_NPS7575__REG_P01_P2_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P01_P2_1_VCA_TOKEN    32'h000000ae
`define NOC2_NPS7575__REG_P01_P2_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P02_P3_0_VCA_TOKEN    32'h000000af
`define NOC2_NPS7575__REG_P02_P3_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P02_P3_1_VCA_TOKEN    32'h000000b0
`define NOC2_NPS7575__REG_P02_P3_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P10_P2_0_VCA_TOKEN    32'h000000b1
`define NOC2_NPS7575__REG_P10_P2_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P10_P2_1_VCA_TOKEN    32'h000000b2
`define NOC2_NPS7575__REG_P10_P2_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P11_P3_0_VCA_TOKEN    32'h000000b3
`define NOC2_NPS7575__REG_P11_P3_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P11_P3_1_VCA_TOKEN    32'h000000b4
`define NOC2_NPS7575__REG_P11_P3_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P12_P0_0_VCA_TOKEN    32'h000000b5
`define NOC2_NPS7575__REG_P12_P0_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P12_P0_1_VCA_TOKEN    32'h000000b6
`define NOC2_NPS7575__REG_P12_P0_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P20_P3_0_VCA_TOKEN    32'h000000b7
`define NOC2_NPS7575__REG_P20_P3_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P20_P3_1_VCA_TOKEN    32'h000000b8
`define NOC2_NPS7575__REG_P20_P3_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P21_P0_0_VCA_TOKEN    32'h000000b9
`define NOC2_NPS7575__REG_P21_P0_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P21_P0_1_VCA_TOKEN    32'h000000ba
`define NOC2_NPS7575__REG_P21_P0_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P22_P1_0_VCA_TOKEN    32'h000000bb
`define NOC2_NPS7575__REG_P22_P1_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P22_P1_1_VCA_TOKEN    32'h000000bc
`define NOC2_NPS7575__REG_P22_P1_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P30_P0_0_VCA_TOKEN    32'h000000bd
`define NOC2_NPS7575__REG_P30_P0_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P30_P0_1_VCA_TOKEN    32'h000000be
`define NOC2_NPS7575__REG_P30_P0_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P31_P1_0_VCA_TOKEN    32'h000000bf
`define NOC2_NPS7575__REG_P31_P1_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P31_P1_1_VCA_TOKEN    32'h000000c0
`define NOC2_NPS7575__REG_P31_P1_1_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P32_P2_0_VCA_TOKEN    32'h000000c1
`define NOC2_NPS7575__REG_P32_P2_0_VCA_TOKEN_SZ 32

`define NOC2_NPS7575__REG_P32_P2_1_VCA_TOKEN    32'h000000c2
`define NOC2_NPS7575__REG_P32_P2_1_VCA_TOKEN_SZ 32

`endif  // B_NOC2_NPS7575_DEFINES_VH