// BLH dynamic attribute configuration look-up table addresses
//

`ifdef B_GTYE5_QUAD_DEFINES_VH
`else
`define B_GTYE5_QUAD_DEFINES_VH

// Look-up table parameters
//

`define GTYE5_QUAD_ADDR_N  792
`define GTYE5_QUAD_ADDR_SZ 32
`define GTYE5_QUAD_DATA_SZ 192

// Attribute addresses
//

`define GTYE5_QUAD__A_CFG0    32'h00000000
`define GTYE5_QUAD__A_CFG0_SZ 32

`define GTYE5_QUAD__A_CFG1    32'h00000001
`define GTYE5_QUAD__A_CFG1_SZ 32

`define GTYE5_QUAD__A_CFG2    32'h00000002
`define GTYE5_QUAD__A_CFG2_SZ 32

`define GTYE5_QUAD__A_CFG3    32'h00000003
`define GTYE5_QUAD__A_CFG3_SZ 32

`define GTYE5_QUAD__A_CFG4    32'h00000004
`define GTYE5_QUAD__A_CFG4_SZ 32

`define GTYE5_QUAD__A_CFG5    32'h00000005
`define GTYE5_QUAD__A_CFG5_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_APT_CFG    32'h00000006
`define GTYE5_QUAD__CH0_ADAPT_APT_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_CAL_CFG    32'h00000007
`define GTYE5_QUAD__CH0_ADAPT_CAL_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_DFE_CFG    32'h00000008
`define GTYE5_QUAD__CH0_ADAPT_DFE_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GC_CFG0    32'h00000009
`define GTYE5_QUAD__CH0_ADAPT_GC_CFG0_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GC_CFG1    32'h0000000a
`define GTYE5_QUAD__CH0_ADAPT_GC_CFG1_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GC_CFG2    32'h0000000b
`define GTYE5_QUAD__CH0_ADAPT_GC_CFG2_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GC_CFG3    32'h0000000c
`define GTYE5_QUAD__CH0_ADAPT_GC_CFG3_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG0    32'h0000000d
`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG0_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG1    32'h0000000e
`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG1_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG2    32'h0000000f
`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG2_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG3    32'h00000010
`define GTYE5_QUAD__CH0_ADAPT_GEN_CFG3_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_H01_CFG    32'h00000011
`define GTYE5_QUAD__CH0_ADAPT_H01_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_H23_CFG    32'h00000012
`define GTYE5_QUAD__CH0_ADAPT_H23_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_H45_CFG    32'h00000013
`define GTYE5_QUAD__CH0_ADAPT_H45_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_H67_CFG    32'h00000014
`define GTYE5_QUAD__CH0_ADAPT_H67_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_H89_CFG    32'h00000015
`define GTYE5_QUAD__CH0_ADAPT_H89_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_HAB_CFG    32'h00000016
`define GTYE5_QUAD__CH0_ADAPT_HAB_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_HCD_CFG    32'h00000017
`define GTYE5_QUAD__CH0_ADAPT_HCD_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_HEF_CFG    32'h00000018
`define GTYE5_QUAD__CH0_ADAPT_HEF_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG0    32'h00000019
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG0_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG1    32'h0000001a
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG1_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG2    32'h0000001b
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG2_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG3    32'h0000001c
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG3_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG4    32'h0000001d
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG4_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KH_CFG5    32'h0000001e
`define GTYE5_QUAD__CH0_ADAPT_KH_CFG5_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KL_CFG0    32'h0000001f
`define GTYE5_QUAD__CH0_ADAPT_KL_CFG0_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_KL_CFG1    32'h00000020
`define GTYE5_QUAD__CH0_ADAPT_KL_CFG1_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG0    32'h00000021
`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG0_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG1    32'h00000022
`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG1_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG2    32'h00000023
`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG2_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG3    32'h00000024
`define GTYE5_QUAD__CH0_ADAPT_LCK_CFG3_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_LOP_CFG    32'h00000025
`define GTYE5_QUAD__CH0_ADAPT_LOP_CFG_SZ 32

`define GTYE5_QUAD__CH0_ADAPT_OS_CFG    32'h00000026
`define GTYE5_QUAD__CH0_ADAPT_OS_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_ILO_CFG    32'h00000027
`define GTYE5_QUAD__CH0_CHCLK_ILO_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_MISC_CFG    32'h00000028
`define GTYE5_QUAD__CH0_CHCLK_MISC_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_RSV_CFG    32'h00000029
`define GTYE5_QUAD__CH0_CHCLK_RSV_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG    32'h0000002a
`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG1    32'h0000002b
`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG1_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG2    32'h0000002c
`define GTYE5_QUAD__CH0_CHCLK_RXCAL_CFG2_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_RXPI_CFG    32'h0000002d
`define GTYE5_QUAD__CH0_CHCLK_RXPI_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_TXCAL_CFG    32'h0000002e
`define GTYE5_QUAD__CH0_CHCLK_TXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH0_CHCLK_TXPI_CFG0    32'h0000002f
`define GTYE5_QUAD__CH0_CHCLK_TXPI_CFG0_SZ 32

`define GTYE5_QUAD__CH0_CHL_RSV_CFG0    32'h00000030
`define GTYE5_QUAD__CH0_CHL_RSV_CFG0_SZ 32

`define GTYE5_QUAD__CH0_CHL_RSV_CFG1    32'h00000031
`define GTYE5_QUAD__CH0_CHL_RSV_CFG1_SZ 32

`define GTYE5_QUAD__CH0_CHL_RSV_CFG2    32'h00000032
`define GTYE5_QUAD__CH0_CHL_RSV_CFG2_SZ 32

`define GTYE5_QUAD__CH0_CHL_RSV_CFG3    32'h00000033
`define GTYE5_QUAD__CH0_CHL_RSV_CFG3_SZ 32

`define GTYE5_QUAD__CH0_CHL_RSV_CFG4    32'h00000034
`define GTYE5_QUAD__CH0_CHL_RSV_CFG4_SZ 32

`define GTYE5_QUAD__CH0_DA_CFG    32'h00000035
`define GTYE5_QUAD__CH0_DA_CFG_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG0    32'h00000036
`define GTYE5_QUAD__CH0_EYESCAN_CFG0_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG1    32'h00000037
`define GTYE5_QUAD__CH0_EYESCAN_CFG1_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG10    32'h00000038
`define GTYE5_QUAD__CH0_EYESCAN_CFG10_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG11    32'h00000039
`define GTYE5_QUAD__CH0_EYESCAN_CFG11_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG12    32'h0000003a
`define GTYE5_QUAD__CH0_EYESCAN_CFG12_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG13    32'h0000003b
`define GTYE5_QUAD__CH0_EYESCAN_CFG13_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG14    32'h0000003c
`define GTYE5_QUAD__CH0_EYESCAN_CFG14_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG15    32'h0000003d
`define GTYE5_QUAD__CH0_EYESCAN_CFG15_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG16    32'h0000003e
`define GTYE5_QUAD__CH0_EYESCAN_CFG16_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG2    32'h0000003f
`define GTYE5_QUAD__CH0_EYESCAN_CFG2_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG3    32'h00000040
`define GTYE5_QUAD__CH0_EYESCAN_CFG3_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG4    32'h00000041
`define GTYE5_QUAD__CH0_EYESCAN_CFG4_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG5    32'h00000042
`define GTYE5_QUAD__CH0_EYESCAN_CFG5_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG6    32'h00000043
`define GTYE5_QUAD__CH0_EYESCAN_CFG6_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG7    32'h00000044
`define GTYE5_QUAD__CH0_EYESCAN_CFG7_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG8    32'h00000045
`define GTYE5_QUAD__CH0_EYESCAN_CFG8_SZ 32

`define GTYE5_QUAD__CH0_EYESCAN_CFG9    32'h00000046
`define GTYE5_QUAD__CH0_EYESCAN_CFG9_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG0    32'h00000047
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG0_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG1    32'h00000048
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG1_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG2    32'h00000049
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG2_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG3    32'h0000004a
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG3_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG4    32'h0000004b
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG4_SZ 32

`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG5    32'h0000004c
`define GTYE5_QUAD__CH0_FABRIC_INTF_CFG5_SZ 32

`define GTYE5_QUAD__CH0_INSTANTIATED    32'h0000004d
`define GTYE5_QUAD__CH0_INSTANTIATED_SZ 1

`define GTYE5_QUAD__CH0_MONITOR_CFG    32'h0000004e
`define GTYE5_QUAD__CH0_MONITOR_CFG_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG0    32'h0000004f
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG0_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG1    32'h00000050
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG1_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG10    32'h00000051
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG10_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG2    32'h00000052
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG2_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG3    32'h00000053
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG3_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG4    32'h00000054
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG4_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG5    32'h00000055
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG5_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG6    32'h00000056
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG6_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG7    32'h00000057
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG7_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG8    32'h00000058
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG8_SZ 32

`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG9    32'h00000059
`define GTYE5_QUAD__CH0_PIPE_CTRL_CFG9_SZ 32

`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG0    32'h0000005a
`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG0_SZ 32

`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG1    32'h0000005b
`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG1_SZ 32

`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG2    32'h0000005c
`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG2_SZ 32

`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG3    32'h0000005d
`define GTYE5_QUAD__CH0_PIPE_TX_EQ_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RESET_BYP_HDSHK_CFG    32'h0000005e
`define GTYE5_QUAD__CH0_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYE5_QUAD__CH0_RESET_CFG    32'h0000005f
`define GTYE5_QUAD__CH0_RESET_CFG_SZ 32

`define GTYE5_QUAD__CH0_RESET_LOOPER_ID_CFG    32'h00000060
`define GTYE5_QUAD__CH0_RESET_LOOPER_ID_CFG_SZ 32

`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG0    32'h00000061
`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG1    32'h00000062
`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG2    32'h00000063
`define GTYE5_QUAD__CH0_RESET_LOOP_ID_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RESET_TIME_CFG0    32'h00000064
`define GTYE5_QUAD__CH0_RESET_TIME_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RESET_TIME_CFG1    32'h00000065
`define GTYE5_QUAD__CH0_RESET_TIME_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RESET_TIME_CFG2    32'h00000066
`define GTYE5_QUAD__CH0_RESET_TIME_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RESET_TIME_CFG3    32'h00000067
`define GTYE5_QUAD__CH0_RESET_TIME_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RXOUTCLK_FREQ    32'h00000068
`define GTYE5_QUAD__CH0_RXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH0_RXOUTCLK_REF_FREQ    32'h00000069
`define GTYE5_QUAD__CH0_RXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH0_RXOUTCLK_REF_SOURCE    32'h0000006a
`define GTYE5_QUAD__CH0_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH0_RX_CDR_CFG0    32'h0000006b
`define GTYE5_QUAD__CH0_RX_CDR_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_CDR_CFG1    32'h0000006c
`define GTYE5_QUAD__CH0_RX_CDR_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_CDR_CFG2    32'h0000006d
`define GTYE5_QUAD__CH0_RX_CDR_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RX_CDR_CFG3    32'h0000006e
`define GTYE5_QUAD__CH0_RX_CDR_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RX_CDR_CFG4    32'h0000006f
`define GTYE5_QUAD__CH0_RX_CDR_CFG4_SZ 32

`define GTYE5_QUAD__CH0_RX_CRC_CFG0    32'h00000070
`define GTYE5_QUAD__CH0_RX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_CRC_CFG1    32'h00000071
`define GTYE5_QUAD__CH0_RX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_CRC_CFG2    32'h00000072
`define GTYE5_QUAD__CH0_RX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RX_CRC_CFG3    32'h00000073
`define GTYE5_QUAD__CH0_RX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RX_CTLE_CFG0    32'h00000074
`define GTYE5_QUAD__CH0_RX_CTLE_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_CTLE_CFG1    32'h00000075
`define GTYE5_QUAD__CH0_RX_CTLE_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_DACI2V_CFG0    32'h00000076
`define GTYE5_QUAD__CH0_RX_DACI2V_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_DATA_RATE    32'h00000077
`define GTYE5_QUAD__CH0_RX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH0_RX_DFE_CFG0    32'h00000078
`define GTYE5_QUAD__CH0_RX_DFE_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG0    32'h00000079
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG1    32'h0000007a
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG2    32'h0000007b
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG3    32'h0000007c
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG4    32'h0000007d
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG5    32'h0000007e
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG6    32'h0000007f
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG7    32'h00000080
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG8    32'h00000081
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG9    32'h00000082
`define GTYE5_QUAD__CH0_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYE5_QUAD__CH0_RX_MISC_CFG0    32'h00000083
`define GTYE5_QUAD__CH0_RX_MISC_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_OOB_CFG0    32'h00000084
`define GTYE5_QUAD__CH0_RX_OOB_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_OOB_CFG1    32'h00000085
`define GTYE5_QUAD__CH0_RX_OOB_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_PAD_CFG0    32'h00000086
`define GTYE5_QUAD__CH0_RX_PAD_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_PAD_CFG1    32'h00000087
`define GTYE5_QUAD__CH0_RX_PAD_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_PCS_CFG0    32'h00000088
`define GTYE5_QUAD__CH0_RX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_PCS_CFG1    32'h00000089
`define GTYE5_QUAD__CH0_RX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_PCS_CFG2    32'h0000008a
`define GTYE5_QUAD__CH0_RX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RX_PCS_CFG3    32'h0000008b
`define GTYE5_QUAD__CH0_RX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RX_PCS_CFG4    32'h0000008c
`define GTYE5_QUAD__CH0_RX_PCS_CFG4_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG0    32'h0000008d
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG1    32'h0000008e
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG2    32'h0000008f
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG3    32'h00000090
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG4    32'h00000091
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG5    32'h00000092
`define GTYE5_QUAD__CH0_RX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH0_SIM_MODE    32'h00000093
`define GTYE5_QUAD__CH0_SIM_MODE_SZ 48

`define GTYE5_QUAD__CH0_SIM_RECEIVER_DETECT_PASS    32'h00000094
`define GTYE5_QUAD__CH0_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYE5_QUAD__CH0_SIM_RESET_SPEEDUP    32'h00000095
`define GTYE5_QUAD__CH0_SIM_RESET_SPEEDUP_SZ 40

`define GTYE5_QUAD__CH0_SIM_TX_EIDLE_DRIVE_LEVEL    32'h00000096
`define GTYE5_QUAD__CH0_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYE5_QUAD__CH0_TXOUTCLK_FREQ    32'h00000097
`define GTYE5_QUAD__CH0_TXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH0_TXOUTCLK_REF_FREQ    32'h00000098
`define GTYE5_QUAD__CH0_TXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH0_TXOUTCLK_REF_SOURCE    32'h00000099
`define GTYE5_QUAD__CH0_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH0_TX_10G_CFG0    32'h0000009a
`define GTYE5_QUAD__CH0_TX_10G_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_10G_CFG1    32'h0000009b
`define GTYE5_QUAD__CH0_TX_10G_CFG1_SZ 32

`define GTYE5_QUAD__CH0_TX_10G_CFG2    32'h0000009c
`define GTYE5_QUAD__CH0_TX_10G_CFG2_SZ 32

`define GTYE5_QUAD__CH0_TX_10G_CFG3    32'h0000009d
`define GTYE5_QUAD__CH0_TX_10G_CFG3_SZ 32

`define GTYE5_QUAD__CH0_TX_ANA_CFG0    32'h0000009e
`define GTYE5_QUAD__CH0_TX_ANA_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_CRC_CFG0    32'h0000009f
`define GTYE5_QUAD__CH0_TX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_CRC_CFG1    32'h000000a0
`define GTYE5_QUAD__CH0_TX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH0_TX_CRC_CFG2    32'h000000a1
`define GTYE5_QUAD__CH0_TX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH0_TX_CRC_CFG3    32'h000000a2
`define GTYE5_QUAD__CH0_TX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH0_TX_DATA_RATE    32'h000000a3
`define GTYE5_QUAD__CH0_TX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH0_TX_DRV_CFG0    32'h000000a4
`define GTYE5_QUAD__CH0_TX_DRV_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_DRV_CFG1    32'h000000a5
`define GTYE5_QUAD__CH0_TX_DRV_CFG1_SZ 32

`define GTYE5_QUAD__CH0_TX_PCS_CFG0    32'h000000a6
`define GTYE5_QUAD__CH0_TX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_PCS_CFG1    32'h000000a7
`define GTYE5_QUAD__CH0_TX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH0_TX_PCS_CFG2    32'h000000a8
`define GTYE5_QUAD__CH0_TX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH0_TX_PCS_CFG3    32'h000000a9
`define GTYE5_QUAD__CH0_TX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG0    32'h000000aa
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG1    32'h000000ab
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG2    32'h000000ac
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG3    32'h000000ad
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG4    32'h000000ae
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG5    32'h000000af
`define GTYE5_QUAD__CH0_TX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH0_TX_PIPPM_CFG    32'h000000b0
`define GTYE5_QUAD__CH0_TX_PIPPM_CFG_SZ 32

`define GTYE5_QUAD__CH0_TX_SER_CFG0    32'h000000b1
`define GTYE5_QUAD__CH0_TX_SER_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_APT_CFG    32'h000000b2
`define GTYE5_QUAD__CH1_ADAPT_APT_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_CAL_CFG    32'h000000b3
`define GTYE5_QUAD__CH1_ADAPT_CAL_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_DFE_CFG    32'h000000b4
`define GTYE5_QUAD__CH1_ADAPT_DFE_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GC_CFG0    32'h000000b5
`define GTYE5_QUAD__CH1_ADAPT_GC_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GC_CFG1    32'h000000b6
`define GTYE5_QUAD__CH1_ADAPT_GC_CFG1_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GC_CFG2    32'h000000b7
`define GTYE5_QUAD__CH1_ADAPT_GC_CFG2_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GC_CFG3    32'h000000b8
`define GTYE5_QUAD__CH1_ADAPT_GC_CFG3_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG0    32'h000000b9
`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG1    32'h000000ba
`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG1_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG2    32'h000000bb
`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG2_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG3    32'h000000bc
`define GTYE5_QUAD__CH1_ADAPT_GEN_CFG3_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_H01_CFG    32'h000000bd
`define GTYE5_QUAD__CH1_ADAPT_H01_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_H23_CFG    32'h000000be
`define GTYE5_QUAD__CH1_ADAPT_H23_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_H45_CFG    32'h000000bf
`define GTYE5_QUAD__CH1_ADAPT_H45_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_H67_CFG    32'h000000c0
`define GTYE5_QUAD__CH1_ADAPT_H67_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_H89_CFG    32'h000000c1
`define GTYE5_QUAD__CH1_ADAPT_H89_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_HAB_CFG    32'h000000c2
`define GTYE5_QUAD__CH1_ADAPT_HAB_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_HCD_CFG    32'h000000c3
`define GTYE5_QUAD__CH1_ADAPT_HCD_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_HEF_CFG    32'h000000c4
`define GTYE5_QUAD__CH1_ADAPT_HEF_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG0    32'h000000c5
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG1    32'h000000c6
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG1_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG2    32'h000000c7
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG2_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG3    32'h000000c8
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG3_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG4    32'h000000c9
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG4_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KH_CFG5    32'h000000ca
`define GTYE5_QUAD__CH1_ADAPT_KH_CFG5_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KL_CFG0    32'h000000cb
`define GTYE5_QUAD__CH1_ADAPT_KL_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_KL_CFG1    32'h000000cc
`define GTYE5_QUAD__CH1_ADAPT_KL_CFG1_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG0    32'h000000cd
`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG0_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG1    32'h000000ce
`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG1_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG2    32'h000000cf
`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG2_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG3    32'h000000d0
`define GTYE5_QUAD__CH1_ADAPT_LCK_CFG3_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_LOP_CFG    32'h000000d1
`define GTYE5_QUAD__CH1_ADAPT_LOP_CFG_SZ 32

`define GTYE5_QUAD__CH1_ADAPT_OS_CFG    32'h000000d2
`define GTYE5_QUAD__CH1_ADAPT_OS_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_ILO_CFG    32'h000000d3
`define GTYE5_QUAD__CH1_CHCLK_ILO_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_MISC_CFG    32'h000000d4
`define GTYE5_QUAD__CH1_CHCLK_MISC_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_RSV_CFG    32'h000000d5
`define GTYE5_QUAD__CH1_CHCLK_RSV_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG    32'h000000d6
`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG1    32'h000000d7
`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG1_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG2    32'h000000d8
`define GTYE5_QUAD__CH1_CHCLK_RXCAL_CFG2_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_RXPI_CFG    32'h000000d9
`define GTYE5_QUAD__CH1_CHCLK_RXPI_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_TXCAL_CFG    32'h000000da
`define GTYE5_QUAD__CH1_CHCLK_TXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH1_CHCLK_TXPI_CFG0    32'h000000db
`define GTYE5_QUAD__CH1_CHCLK_TXPI_CFG0_SZ 32

`define GTYE5_QUAD__CH1_CHL_RSV_CFG0    32'h000000dc
`define GTYE5_QUAD__CH1_CHL_RSV_CFG0_SZ 32

`define GTYE5_QUAD__CH1_CHL_RSV_CFG1    32'h000000dd
`define GTYE5_QUAD__CH1_CHL_RSV_CFG1_SZ 32

`define GTYE5_QUAD__CH1_CHL_RSV_CFG2    32'h000000de
`define GTYE5_QUAD__CH1_CHL_RSV_CFG2_SZ 32

`define GTYE5_QUAD__CH1_CHL_RSV_CFG3    32'h000000df
`define GTYE5_QUAD__CH1_CHL_RSV_CFG3_SZ 32

`define GTYE5_QUAD__CH1_CHL_RSV_CFG4    32'h000000e0
`define GTYE5_QUAD__CH1_CHL_RSV_CFG4_SZ 32

`define GTYE5_QUAD__CH1_DA_CFG    32'h000000e1
`define GTYE5_QUAD__CH1_DA_CFG_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG0    32'h000000e2
`define GTYE5_QUAD__CH1_EYESCAN_CFG0_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG1    32'h000000e3
`define GTYE5_QUAD__CH1_EYESCAN_CFG1_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG10    32'h000000e4
`define GTYE5_QUAD__CH1_EYESCAN_CFG10_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG11    32'h000000e5
`define GTYE5_QUAD__CH1_EYESCAN_CFG11_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG12    32'h000000e6
`define GTYE5_QUAD__CH1_EYESCAN_CFG12_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG13    32'h000000e7
`define GTYE5_QUAD__CH1_EYESCAN_CFG13_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG14    32'h000000e8
`define GTYE5_QUAD__CH1_EYESCAN_CFG14_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG15    32'h000000e9
`define GTYE5_QUAD__CH1_EYESCAN_CFG15_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG16    32'h000000ea
`define GTYE5_QUAD__CH1_EYESCAN_CFG16_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG2    32'h000000eb
`define GTYE5_QUAD__CH1_EYESCAN_CFG2_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG3    32'h000000ec
`define GTYE5_QUAD__CH1_EYESCAN_CFG3_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG4    32'h000000ed
`define GTYE5_QUAD__CH1_EYESCAN_CFG4_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG5    32'h000000ee
`define GTYE5_QUAD__CH1_EYESCAN_CFG5_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG6    32'h000000ef
`define GTYE5_QUAD__CH1_EYESCAN_CFG6_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG7    32'h000000f0
`define GTYE5_QUAD__CH1_EYESCAN_CFG7_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG8    32'h000000f1
`define GTYE5_QUAD__CH1_EYESCAN_CFG8_SZ 32

`define GTYE5_QUAD__CH1_EYESCAN_CFG9    32'h000000f2
`define GTYE5_QUAD__CH1_EYESCAN_CFG9_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG0    32'h000000f3
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG0_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG1    32'h000000f4
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG1_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG2    32'h000000f5
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG2_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG3    32'h000000f6
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG3_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG4    32'h000000f7
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG4_SZ 32

`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG5    32'h000000f8
`define GTYE5_QUAD__CH1_FABRIC_INTF_CFG5_SZ 32

`define GTYE5_QUAD__CH1_INSTANTIATED    32'h000000f9
`define GTYE5_QUAD__CH1_INSTANTIATED_SZ 1

`define GTYE5_QUAD__CH1_MONITOR_CFG    32'h000000fa
`define GTYE5_QUAD__CH1_MONITOR_CFG_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG0    32'h000000fb
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG0_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG1    32'h000000fc
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG1_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG10    32'h000000fd
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG10_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG2    32'h000000fe
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG2_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG3    32'h000000ff
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG3_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG4    32'h00000100
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG4_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG5    32'h00000101
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG5_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG6    32'h00000102
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG6_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG7    32'h00000103
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG7_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG8    32'h00000104
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG8_SZ 32

`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG9    32'h00000105
`define GTYE5_QUAD__CH1_PIPE_CTRL_CFG9_SZ 32

`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG0    32'h00000106
`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG0_SZ 32

`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG1    32'h00000107
`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG1_SZ 32

`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG2    32'h00000108
`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG2_SZ 32

`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG3    32'h00000109
`define GTYE5_QUAD__CH1_PIPE_TX_EQ_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RESET_BYP_HDSHK_CFG    32'h0000010a
`define GTYE5_QUAD__CH1_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYE5_QUAD__CH1_RESET_CFG    32'h0000010b
`define GTYE5_QUAD__CH1_RESET_CFG_SZ 32

`define GTYE5_QUAD__CH1_RESET_LOOPER_ID_CFG    32'h0000010c
`define GTYE5_QUAD__CH1_RESET_LOOPER_ID_CFG_SZ 32

`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG0    32'h0000010d
`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG1    32'h0000010e
`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG2    32'h0000010f
`define GTYE5_QUAD__CH1_RESET_LOOP_ID_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RESET_TIME_CFG0    32'h00000110
`define GTYE5_QUAD__CH1_RESET_TIME_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RESET_TIME_CFG1    32'h00000111
`define GTYE5_QUAD__CH1_RESET_TIME_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RESET_TIME_CFG2    32'h00000112
`define GTYE5_QUAD__CH1_RESET_TIME_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RESET_TIME_CFG3    32'h00000113
`define GTYE5_QUAD__CH1_RESET_TIME_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RXOUTCLK_FREQ    32'h00000114
`define GTYE5_QUAD__CH1_RXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH1_RXOUTCLK_REF_FREQ    32'h00000115
`define GTYE5_QUAD__CH1_RXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH1_RXOUTCLK_REF_SOURCE    32'h00000116
`define GTYE5_QUAD__CH1_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH1_RX_CDR_CFG0    32'h00000117
`define GTYE5_QUAD__CH1_RX_CDR_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_CDR_CFG1    32'h00000118
`define GTYE5_QUAD__CH1_RX_CDR_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_CDR_CFG2    32'h00000119
`define GTYE5_QUAD__CH1_RX_CDR_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RX_CDR_CFG3    32'h0000011a
`define GTYE5_QUAD__CH1_RX_CDR_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RX_CDR_CFG4    32'h0000011b
`define GTYE5_QUAD__CH1_RX_CDR_CFG4_SZ 32

`define GTYE5_QUAD__CH1_RX_CRC_CFG0    32'h0000011c
`define GTYE5_QUAD__CH1_RX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_CRC_CFG1    32'h0000011d
`define GTYE5_QUAD__CH1_RX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_CRC_CFG2    32'h0000011e
`define GTYE5_QUAD__CH1_RX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RX_CRC_CFG3    32'h0000011f
`define GTYE5_QUAD__CH1_RX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RX_CTLE_CFG0    32'h00000120
`define GTYE5_QUAD__CH1_RX_CTLE_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_CTLE_CFG1    32'h00000121
`define GTYE5_QUAD__CH1_RX_CTLE_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_DACI2V_CFG0    32'h00000122
`define GTYE5_QUAD__CH1_RX_DACI2V_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_DATA_RATE    32'h00000123
`define GTYE5_QUAD__CH1_RX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH1_RX_DFE_CFG0    32'h00000124
`define GTYE5_QUAD__CH1_RX_DFE_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG0    32'h00000125
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG1    32'h00000126
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG2    32'h00000127
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG3    32'h00000128
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG4    32'h00000129
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG5    32'h0000012a
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG6    32'h0000012b
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG7    32'h0000012c
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG8    32'h0000012d
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG9    32'h0000012e
`define GTYE5_QUAD__CH1_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYE5_QUAD__CH1_RX_MISC_CFG0    32'h0000012f
`define GTYE5_QUAD__CH1_RX_MISC_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_OOB_CFG0    32'h00000130
`define GTYE5_QUAD__CH1_RX_OOB_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_OOB_CFG1    32'h00000131
`define GTYE5_QUAD__CH1_RX_OOB_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_PAD_CFG0    32'h00000132
`define GTYE5_QUAD__CH1_RX_PAD_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_PAD_CFG1    32'h00000133
`define GTYE5_QUAD__CH1_RX_PAD_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_PCS_CFG0    32'h00000134
`define GTYE5_QUAD__CH1_RX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_PCS_CFG1    32'h00000135
`define GTYE5_QUAD__CH1_RX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_PCS_CFG2    32'h00000136
`define GTYE5_QUAD__CH1_RX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RX_PCS_CFG3    32'h00000137
`define GTYE5_QUAD__CH1_RX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RX_PCS_CFG4    32'h00000138
`define GTYE5_QUAD__CH1_RX_PCS_CFG4_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG0    32'h00000139
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG1    32'h0000013a
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG2    32'h0000013b
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG3    32'h0000013c
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG4    32'h0000013d
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG5    32'h0000013e
`define GTYE5_QUAD__CH1_RX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH1_SIM_MODE    32'h0000013f
`define GTYE5_QUAD__CH1_SIM_MODE_SZ 48

`define GTYE5_QUAD__CH1_SIM_RECEIVER_DETECT_PASS    32'h00000140
`define GTYE5_QUAD__CH1_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYE5_QUAD__CH1_SIM_RESET_SPEEDUP    32'h00000141
`define GTYE5_QUAD__CH1_SIM_RESET_SPEEDUP_SZ 40

`define GTYE5_QUAD__CH1_SIM_TX_EIDLE_DRIVE_LEVEL    32'h00000142
`define GTYE5_QUAD__CH1_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYE5_QUAD__CH1_TXOUTCLK_FREQ    32'h00000143
`define GTYE5_QUAD__CH1_TXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH1_TXOUTCLK_REF_FREQ    32'h00000144
`define GTYE5_QUAD__CH1_TXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH1_TXOUTCLK_REF_SOURCE    32'h00000145
`define GTYE5_QUAD__CH1_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH1_TX_10G_CFG0    32'h00000146
`define GTYE5_QUAD__CH1_TX_10G_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_10G_CFG1    32'h00000147
`define GTYE5_QUAD__CH1_TX_10G_CFG1_SZ 32

`define GTYE5_QUAD__CH1_TX_10G_CFG2    32'h00000148
`define GTYE5_QUAD__CH1_TX_10G_CFG2_SZ 32

`define GTYE5_QUAD__CH1_TX_10G_CFG3    32'h00000149
`define GTYE5_QUAD__CH1_TX_10G_CFG3_SZ 32

`define GTYE5_QUAD__CH1_TX_ANA_CFG0    32'h0000014a
`define GTYE5_QUAD__CH1_TX_ANA_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_CRC_CFG0    32'h0000014b
`define GTYE5_QUAD__CH1_TX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_CRC_CFG1    32'h0000014c
`define GTYE5_QUAD__CH1_TX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH1_TX_CRC_CFG2    32'h0000014d
`define GTYE5_QUAD__CH1_TX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH1_TX_CRC_CFG3    32'h0000014e
`define GTYE5_QUAD__CH1_TX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH1_TX_DATA_RATE    32'h0000014f
`define GTYE5_QUAD__CH1_TX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH1_TX_DRV_CFG0    32'h00000150
`define GTYE5_QUAD__CH1_TX_DRV_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_DRV_CFG1    32'h00000151
`define GTYE5_QUAD__CH1_TX_DRV_CFG1_SZ 32

`define GTYE5_QUAD__CH1_TX_PCS_CFG0    32'h00000152
`define GTYE5_QUAD__CH1_TX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_PCS_CFG1    32'h00000153
`define GTYE5_QUAD__CH1_TX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH1_TX_PCS_CFG2    32'h00000154
`define GTYE5_QUAD__CH1_TX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH1_TX_PCS_CFG3    32'h00000155
`define GTYE5_QUAD__CH1_TX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG0    32'h00000156
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG1    32'h00000157
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG2    32'h00000158
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG3    32'h00000159
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG4    32'h0000015a
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG5    32'h0000015b
`define GTYE5_QUAD__CH1_TX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH1_TX_PIPPM_CFG    32'h0000015c
`define GTYE5_QUAD__CH1_TX_PIPPM_CFG_SZ 32

`define GTYE5_QUAD__CH1_TX_SER_CFG0    32'h0000015d
`define GTYE5_QUAD__CH1_TX_SER_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_APT_CFG    32'h0000015e
`define GTYE5_QUAD__CH2_ADAPT_APT_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_CAL_CFG    32'h0000015f
`define GTYE5_QUAD__CH2_ADAPT_CAL_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_DFE_CFG    32'h00000160
`define GTYE5_QUAD__CH2_ADAPT_DFE_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GC_CFG0    32'h00000161
`define GTYE5_QUAD__CH2_ADAPT_GC_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GC_CFG1    32'h00000162
`define GTYE5_QUAD__CH2_ADAPT_GC_CFG1_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GC_CFG2    32'h00000163
`define GTYE5_QUAD__CH2_ADAPT_GC_CFG2_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GC_CFG3    32'h00000164
`define GTYE5_QUAD__CH2_ADAPT_GC_CFG3_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG0    32'h00000165
`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG1    32'h00000166
`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG1_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG2    32'h00000167
`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG2_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG3    32'h00000168
`define GTYE5_QUAD__CH2_ADAPT_GEN_CFG3_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_H01_CFG    32'h00000169
`define GTYE5_QUAD__CH2_ADAPT_H01_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_H23_CFG    32'h0000016a
`define GTYE5_QUAD__CH2_ADAPT_H23_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_H45_CFG    32'h0000016b
`define GTYE5_QUAD__CH2_ADAPT_H45_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_H67_CFG    32'h0000016c
`define GTYE5_QUAD__CH2_ADAPT_H67_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_H89_CFG    32'h0000016d
`define GTYE5_QUAD__CH2_ADAPT_H89_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_HAB_CFG    32'h0000016e
`define GTYE5_QUAD__CH2_ADAPT_HAB_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_HCD_CFG    32'h0000016f
`define GTYE5_QUAD__CH2_ADAPT_HCD_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_HEF_CFG    32'h00000170
`define GTYE5_QUAD__CH2_ADAPT_HEF_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG0    32'h00000171
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG1    32'h00000172
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG1_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG2    32'h00000173
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG2_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG3    32'h00000174
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG3_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG4    32'h00000175
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG4_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KH_CFG5    32'h00000176
`define GTYE5_QUAD__CH2_ADAPT_KH_CFG5_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KL_CFG0    32'h00000177
`define GTYE5_QUAD__CH2_ADAPT_KL_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_KL_CFG1    32'h00000178
`define GTYE5_QUAD__CH2_ADAPT_KL_CFG1_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG0    32'h00000179
`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG0_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG1    32'h0000017a
`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG1_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG2    32'h0000017b
`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG2_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG3    32'h0000017c
`define GTYE5_QUAD__CH2_ADAPT_LCK_CFG3_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_LOP_CFG    32'h0000017d
`define GTYE5_QUAD__CH2_ADAPT_LOP_CFG_SZ 32

`define GTYE5_QUAD__CH2_ADAPT_OS_CFG    32'h0000017e
`define GTYE5_QUAD__CH2_ADAPT_OS_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_ILO_CFG    32'h0000017f
`define GTYE5_QUAD__CH2_CHCLK_ILO_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_MISC_CFG    32'h00000180
`define GTYE5_QUAD__CH2_CHCLK_MISC_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_RSV_CFG    32'h00000181
`define GTYE5_QUAD__CH2_CHCLK_RSV_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG    32'h00000182
`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG1    32'h00000183
`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG1_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG2    32'h00000184
`define GTYE5_QUAD__CH2_CHCLK_RXCAL_CFG2_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_RXPI_CFG    32'h00000185
`define GTYE5_QUAD__CH2_CHCLK_RXPI_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_TXCAL_CFG    32'h00000186
`define GTYE5_QUAD__CH2_CHCLK_TXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH2_CHCLK_TXPI_CFG0    32'h00000187
`define GTYE5_QUAD__CH2_CHCLK_TXPI_CFG0_SZ 32

`define GTYE5_QUAD__CH2_CHL_RSV_CFG0    32'h00000188
`define GTYE5_QUAD__CH2_CHL_RSV_CFG0_SZ 32

`define GTYE5_QUAD__CH2_CHL_RSV_CFG1    32'h00000189
`define GTYE5_QUAD__CH2_CHL_RSV_CFG1_SZ 32

`define GTYE5_QUAD__CH2_CHL_RSV_CFG2    32'h0000018a
`define GTYE5_QUAD__CH2_CHL_RSV_CFG2_SZ 32

`define GTYE5_QUAD__CH2_CHL_RSV_CFG3    32'h0000018b
`define GTYE5_QUAD__CH2_CHL_RSV_CFG3_SZ 32

`define GTYE5_QUAD__CH2_CHL_RSV_CFG4    32'h0000018c
`define GTYE5_QUAD__CH2_CHL_RSV_CFG4_SZ 32

`define GTYE5_QUAD__CH2_DA_CFG    32'h0000018d
`define GTYE5_QUAD__CH2_DA_CFG_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG0    32'h0000018e
`define GTYE5_QUAD__CH2_EYESCAN_CFG0_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG1    32'h0000018f
`define GTYE5_QUAD__CH2_EYESCAN_CFG1_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG10    32'h00000190
`define GTYE5_QUAD__CH2_EYESCAN_CFG10_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG11    32'h00000191
`define GTYE5_QUAD__CH2_EYESCAN_CFG11_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG12    32'h00000192
`define GTYE5_QUAD__CH2_EYESCAN_CFG12_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG13    32'h00000193
`define GTYE5_QUAD__CH2_EYESCAN_CFG13_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG14    32'h00000194
`define GTYE5_QUAD__CH2_EYESCAN_CFG14_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG15    32'h00000195
`define GTYE5_QUAD__CH2_EYESCAN_CFG15_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG16    32'h00000196
`define GTYE5_QUAD__CH2_EYESCAN_CFG16_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG2    32'h00000197
`define GTYE5_QUAD__CH2_EYESCAN_CFG2_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG3    32'h00000198
`define GTYE5_QUAD__CH2_EYESCAN_CFG3_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG4    32'h00000199
`define GTYE5_QUAD__CH2_EYESCAN_CFG4_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG5    32'h0000019a
`define GTYE5_QUAD__CH2_EYESCAN_CFG5_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG6    32'h0000019b
`define GTYE5_QUAD__CH2_EYESCAN_CFG6_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG7    32'h0000019c
`define GTYE5_QUAD__CH2_EYESCAN_CFG7_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG8    32'h0000019d
`define GTYE5_QUAD__CH2_EYESCAN_CFG8_SZ 32

`define GTYE5_QUAD__CH2_EYESCAN_CFG9    32'h0000019e
`define GTYE5_QUAD__CH2_EYESCAN_CFG9_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG0    32'h0000019f
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG0_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG1    32'h000001a0
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG1_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG2    32'h000001a1
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG2_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG3    32'h000001a2
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG3_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG4    32'h000001a3
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG4_SZ 32

`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG5    32'h000001a4
`define GTYE5_QUAD__CH2_FABRIC_INTF_CFG5_SZ 32

`define GTYE5_QUAD__CH2_INSTANTIATED    32'h000001a5
`define GTYE5_QUAD__CH2_INSTANTIATED_SZ 1

`define GTYE5_QUAD__CH2_MONITOR_CFG    32'h000001a6
`define GTYE5_QUAD__CH2_MONITOR_CFG_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG0    32'h000001a7
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG0_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG1    32'h000001a8
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG1_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG10    32'h000001a9
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG10_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG2    32'h000001aa
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG2_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG3    32'h000001ab
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG3_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG4    32'h000001ac
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG4_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG5    32'h000001ad
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG5_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG6    32'h000001ae
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG6_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG7    32'h000001af
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG7_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG8    32'h000001b0
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG8_SZ 32

`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG9    32'h000001b1
`define GTYE5_QUAD__CH2_PIPE_CTRL_CFG9_SZ 32

`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG0    32'h000001b2
`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG0_SZ 32

`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG1    32'h000001b3
`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG1_SZ 32

`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG2    32'h000001b4
`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG2_SZ 32

`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG3    32'h000001b5
`define GTYE5_QUAD__CH2_PIPE_TX_EQ_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RESET_BYP_HDSHK_CFG    32'h000001b6
`define GTYE5_QUAD__CH2_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYE5_QUAD__CH2_RESET_CFG    32'h000001b7
`define GTYE5_QUAD__CH2_RESET_CFG_SZ 32

`define GTYE5_QUAD__CH2_RESET_LOOPER_ID_CFG    32'h000001b8
`define GTYE5_QUAD__CH2_RESET_LOOPER_ID_CFG_SZ 32

`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG0    32'h000001b9
`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG1    32'h000001ba
`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG2    32'h000001bb
`define GTYE5_QUAD__CH2_RESET_LOOP_ID_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RESET_TIME_CFG0    32'h000001bc
`define GTYE5_QUAD__CH2_RESET_TIME_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RESET_TIME_CFG1    32'h000001bd
`define GTYE5_QUAD__CH2_RESET_TIME_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RESET_TIME_CFG2    32'h000001be
`define GTYE5_QUAD__CH2_RESET_TIME_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RESET_TIME_CFG3    32'h000001bf
`define GTYE5_QUAD__CH2_RESET_TIME_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RXOUTCLK_FREQ    32'h000001c0
`define GTYE5_QUAD__CH2_RXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH2_RXOUTCLK_REF_FREQ    32'h000001c1
`define GTYE5_QUAD__CH2_RXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH2_RXOUTCLK_REF_SOURCE    32'h000001c2
`define GTYE5_QUAD__CH2_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH2_RX_CDR_CFG0    32'h000001c3
`define GTYE5_QUAD__CH2_RX_CDR_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_CDR_CFG1    32'h000001c4
`define GTYE5_QUAD__CH2_RX_CDR_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_CDR_CFG2    32'h000001c5
`define GTYE5_QUAD__CH2_RX_CDR_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RX_CDR_CFG3    32'h000001c6
`define GTYE5_QUAD__CH2_RX_CDR_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RX_CDR_CFG4    32'h000001c7
`define GTYE5_QUAD__CH2_RX_CDR_CFG4_SZ 32

`define GTYE5_QUAD__CH2_RX_CRC_CFG0    32'h000001c8
`define GTYE5_QUAD__CH2_RX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_CRC_CFG1    32'h000001c9
`define GTYE5_QUAD__CH2_RX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_CRC_CFG2    32'h000001ca
`define GTYE5_QUAD__CH2_RX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RX_CRC_CFG3    32'h000001cb
`define GTYE5_QUAD__CH2_RX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RX_CTLE_CFG0    32'h000001cc
`define GTYE5_QUAD__CH2_RX_CTLE_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_CTLE_CFG1    32'h000001cd
`define GTYE5_QUAD__CH2_RX_CTLE_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_DACI2V_CFG0    32'h000001ce
`define GTYE5_QUAD__CH2_RX_DACI2V_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_DATA_RATE    32'h000001cf
`define GTYE5_QUAD__CH2_RX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH2_RX_DFE_CFG0    32'h000001d0
`define GTYE5_QUAD__CH2_RX_DFE_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG0    32'h000001d1
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG1    32'h000001d2
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG2    32'h000001d3
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG3    32'h000001d4
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG4    32'h000001d5
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG5    32'h000001d6
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG6    32'h000001d7
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG7    32'h000001d8
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG8    32'h000001d9
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG9    32'h000001da
`define GTYE5_QUAD__CH2_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYE5_QUAD__CH2_RX_MISC_CFG0    32'h000001db
`define GTYE5_QUAD__CH2_RX_MISC_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_OOB_CFG0    32'h000001dc
`define GTYE5_QUAD__CH2_RX_OOB_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_OOB_CFG1    32'h000001dd
`define GTYE5_QUAD__CH2_RX_OOB_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_PAD_CFG0    32'h000001de
`define GTYE5_QUAD__CH2_RX_PAD_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_PAD_CFG1    32'h000001df
`define GTYE5_QUAD__CH2_RX_PAD_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_PCS_CFG0    32'h000001e0
`define GTYE5_QUAD__CH2_RX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_PCS_CFG1    32'h000001e1
`define GTYE5_QUAD__CH2_RX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_PCS_CFG2    32'h000001e2
`define GTYE5_QUAD__CH2_RX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RX_PCS_CFG3    32'h000001e3
`define GTYE5_QUAD__CH2_RX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RX_PCS_CFG4    32'h000001e4
`define GTYE5_QUAD__CH2_RX_PCS_CFG4_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG0    32'h000001e5
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG1    32'h000001e6
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG2    32'h000001e7
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG3    32'h000001e8
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG4    32'h000001e9
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG5    32'h000001ea
`define GTYE5_QUAD__CH2_RX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH2_SIM_MODE    32'h000001eb
`define GTYE5_QUAD__CH2_SIM_MODE_SZ 48

`define GTYE5_QUAD__CH2_SIM_RECEIVER_DETECT_PASS    32'h000001ec
`define GTYE5_QUAD__CH2_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYE5_QUAD__CH2_SIM_RESET_SPEEDUP    32'h000001ed
`define GTYE5_QUAD__CH2_SIM_RESET_SPEEDUP_SZ 40

`define GTYE5_QUAD__CH2_SIM_TX_EIDLE_DRIVE_LEVEL    32'h000001ee
`define GTYE5_QUAD__CH2_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYE5_QUAD__CH2_TXOUTCLK_FREQ    32'h000001ef
`define GTYE5_QUAD__CH2_TXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH2_TXOUTCLK_REF_FREQ    32'h000001f0
`define GTYE5_QUAD__CH2_TXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH2_TXOUTCLK_REF_SOURCE    32'h000001f1
`define GTYE5_QUAD__CH2_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH2_TX_10G_CFG0    32'h000001f2
`define GTYE5_QUAD__CH2_TX_10G_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_10G_CFG1    32'h000001f3
`define GTYE5_QUAD__CH2_TX_10G_CFG1_SZ 32

`define GTYE5_QUAD__CH2_TX_10G_CFG2    32'h000001f4
`define GTYE5_QUAD__CH2_TX_10G_CFG2_SZ 32

`define GTYE5_QUAD__CH2_TX_10G_CFG3    32'h000001f5
`define GTYE5_QUAD__CH2_TX_10G_CFG3_SZ 32

`define GTYE5_QUAD__CH2_TX_ANA_CFG0    32'h000001f6
`define GTYE5_QUAD__CH2_TX_ANA_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_CRC_CFG0    32'h000001f7
`define GTYE5_QUAD__CH2_TX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_CRC_CFG1    32'h000001f8
`define GTYE5_QUAD__CH2_TX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH2_TX_CRC_CFG2    32'h000001f9
`define GTYE5_QUAD__CH2_TX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH2_TX_CRC_CFG3    32'h000001fa
`define GTYE5_QUAD__CH2_TX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH2_TX_DATA_RATE    32'h000001fb
`define GTYE5_QUAD__CH2_TX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH2_TX_DRV_CFG0    32'h000001fc
`define GTYE5_QUAD__CH2_TX_DRV_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_DRV_CFG1    32'h000001fd
`define GTYE5_QUAD__CH2_TX_DRV_CFG1_SZ 32

`define GTYE5_QUAD__CH2_TX_PCS_CFG0    32'h000001fe
`define GTYE5_QUAD__CH2_TX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_PCS_CFG1    32'h000001ff
`define GTYE5_QUAD__CH2_TX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH2_TX_PCS_CFG2    32'h00000200
`define GTYE5_QUAD__CH2_TX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH2_TX_PCS_CFG3    32'h00000201
`define GTYE5_QUAD__CH2_TX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG0    32'h00000202
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG1    32'h00000203
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG2    32'h00000204
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG3    32'h00000205
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG4    32'h00000206
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG5    32'h00000207
`define GTYE5_QUAD__CH2_TX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH2_TX_PIPPM_CFG    32'h00000208
`define GTYE5_QUAD__CH2_TX_PIPPM_CFG_SZ 32

`define GTYE5_QUAD__CH2_TX_SER_CFG0    32'h00000209
`define GTYE5_QUAD__CH2_TX_SER_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_APT_CFG    32'h0000020a
`define GTYE5_QUAD__CH3_ADAPT_APT_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_CAL_CFG    32'h0000020b
`define GTYE5_QUAD__CH3_ADAPT_CAL_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_DFE_CFG    32'h0000020c
`define GTYE5_QUAD__CH3_ADAPT_DFE_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GC_CFG0    32'h0000020d
`define GTYE5_QUAD__CH3_ADAPT_GC_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GC_CFG1    32'h0000020e
`define GTYE5_QUAD__CH3_ADAPT_GC_CFG1_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GC_CFG2    32'h0000020f
`define GTYE5_QUAD__CH3_ADAPT_GC_CFG2_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GC_CFG3    32'h00000210
`define GTYE5_QUAD__CH3_ADAPT_GC_CFG3_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG0    32'h00000211
`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG1    32'h00000212
`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG1_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG2    32'h00000213
`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG2_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG3    32'h00000214
`define GTYE5_QUAD__CH3_ADAPT_GEN_CFG3_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_H01_CFG    32'h00000215
`define GTYE5_QUAD__CH3_ADAPT_H01_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_H23_CFG    32'h00000216
`define GTYE5_QUAD__CH3_ADAPT_H23_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_H45_CFG    32'h00000217
`define GTYE5_QUAD__CH3_ADAPT_H45_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_H67_CFG    32'h00000218
`define GTYE5_QUAD__CH3_ADAPT_H67_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_H89_CFG    32'h00000219
`define GTYE5_QUAD__CH3_ADAPT_H89_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_HAB_CFG    32'h0000021a
`define GTYE5_QUAD__CH3_ADAPT_HAB_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_HCD_CFG    32'h0000021b
`define GTYE5_QUAD__CH3_ADAPT_HCD_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_HEF_CFG    32'h0000021c
`define GTYE5_QUAD__CH3_ADAPT_HEF_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG0    32'h0000021d
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG1    32'h0000021e
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG1_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG2    32'h0000021f
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG2_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG3    32'h00000220
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG3_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG4    32'h00000221
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG4_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KH_CFG5    32'h00000222
`define GTYE5_QUAD__CH3_ADAPT_KH_CFG5_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KL_CFG0    32'h00000223
`define GTYE5_QUAD__CH3_ADAPT_KL_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_KL_CFG1    32'h00000224
`define GTYE5_QUAD__CH3_ADAPT_KL_CFG1_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG0    32'h00000225
`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG0_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG1    32'h00000226
`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG1_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG2    32'h00000227
`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG2_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG3    32'h00000228
`define GTYE5_QUAD__CH3_ADAPT_LCK_CFG3_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_LOP_CFG    32'h00000229
`define GTYE5_QUAD__CH3_ADAPT_LOP_CFG_SZ 32

`define GTYE5_QUAD__CH3_ADAPT_OS_CFG    32'h0000022a
`define GTYE5_QUAD__CH3_ADAPT_OS_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_ILO_CFG    32'h0000022b
`define GTYE5_QUAD__CH3_CHCLK_ILO_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_MISC_CFG    32'h0000022c
`define GTYE5_QUAD__CH3_CHCLK_MISC_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_RSV_CFG    32'h0000022d
`define GTYE5_QUAD__CH3_CHCLK_RSV_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG    32'h0000022e
`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG1    32'h0000022f
`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG1_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG2    32'h00000230
`define GTYE5_QUAD__CH3_CHCLK_RXCAL_CFG2_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_RXPI_CFG    32'h00000231
`define GTYE5_QUAD__CH3_CHCLK_RXPI_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_TXCAL_CFG    32'h00000232
`define GTYE5_QUAD__CH3_CHCLK_TXCAL_CFG_SZ 32

`define GTYE5_QUAD__CH3_CHCLK_TXPI_CFG0    32'h00000233
`define GTYE5_QUAD__CH3_CHCLK_TXPI_CFG0_SZ 32

`define GTYE5_QUAD__CH3_CHL_RSV_CFG0    32'h00000234
`define GTYE5_QUAD__CH3_CHL_RSV_CFG0_SZ 32

`define GTYE5_QUAD__CH3_CHL_RSV_CFG1    32'h00000235
`define GTYE5_QUAD__CH3_CHL_RSV_CFG1_SZ 32

`define GTYE5_QUAD__CH3_CHL_RSV_CFG2    32'h00000236
`define GTYE5_QUAD__CH3_CHL_RSV_CFG2_SZ 32

`define GTYE5_QUAD__CH3_CHL_RSV_CFG3    32'h00000237
`define GTYE5_QUAD__CH3_CHL_RSV_CFG3_SZ 32

`define GTYE5_QUAD__CH3_CHL_RSV_CFG4    32'h00000238
`define GTYE5_QUAD__CH3_CHL_RSV_CFG4_SZ 32

`define GTYE5_QUAD__CH3_DA_CFG    32'h00000239
`define GTYE5_QUAD__CH3_DA_CFG_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG0    32'h0000023a
`define GTYE5_QUAD__CH3_EYESCAN_CFG0_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG1    32'h0000023b
`define GTYE5_QUAD__CH3_EYESCAN_CFG1_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG10    32'h0000023c
`define GTYE5_QUAD__CH3_EYESCAN_CFG10_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG11    32'h0000023d
`define GTYE5_QUAD__CH3_EYESCAN_CFG11_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG12    32'h0000023e
`define GTYE5_QUAD__CH3_EYESCAN_CFG12_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG13    32'h0000023f
`define GTYE5_QUAD__CH3_EYESCAN_CFG13_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG14    32'h00000240
`define GTYE5_QUAD__CH3_EYESCAN_CFG14_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG15    32'h00000241
`define GTYE5_QUAD__CH3_EYESCAN_CFG15_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG16    32'h00000242
`define GTYE5_QUAD__CH3_EYESCAN_CFG16_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG2    32'h00000243
`define GTYE5_QUAD__CH3_EYESCAN_CFG2_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG3    32'h00000244
`define GTYE5_QUAD__CH3_EYESCAN_CFG3_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG4    32'h00000245
`define GTYE5_QUAD__CH3_EYESCAN_CFG4_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG5    32'h00000246
`define GTYE5_QUAD__CH3_EYESCAN_CFG5_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG6    32'h00000247
`define GTYE5_QUAD__CH3_EYESCAN_CFG6_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG7    32'h00000248
`define GTYE5_QUAD__CH3_EYESCAN_CFG7_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG8    32'h00000249
`define GTYE5_QUAD__CH3_EYESCAN_CFG8_SZ 32

`define GTYE5_QUAD__CH3_EYESCAN_CFG9    32'h0000024a
`define GTYE5_QUAD__CH3_EYESCAN_CFG9_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG0    32'h0000024b
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG0_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG1    32'h0000024c
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG1_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG2    32'h0000024d
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG2_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG3    32'h0000024e
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG3_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG4    32'h0000024f
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG4_SZ 32

`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG5    32'h00000250
`define GTYE5_QUAD__CH3_FABRIC_INTF_CFG5_SZ 32

`define GTYE5_QUAD__CH3_INSTANTIATED    32'h00000251
`define GTYE5_QUAD__CH3_INSTANTIATED_SZ 1

`define GTYE5_QUAD__CH3_MONITOR_CFG    32'h00000252
`define GTYE5_QUAD__CH3_MONITOR_CFG_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG0    32'h00000253
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG0_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG1    32'h00000254
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG1_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG10    32'h00000255
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG10_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG2    32'h00000256
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG2_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG3    32'h00000257
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG3_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG4    32'h00000258
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG4_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG5    32'h00000259
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG5_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG6    32'h0000025a
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG6_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG7    32'h0000025b
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG7_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG8    32'h0000025c
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG8_SZ 32

`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG9    32'h0000025d
`define GTYE5_QUAD__CH3_PIPE_CTRL_CFG9_SZ 32

`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG0    32'h0000025e
`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG0_SZ 32

`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG1    32'h0000025f
`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG1_SZ 32

`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG2    32'h00000260
`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG2_SZ 32

`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG3    32'h00000261
`define GTYE5_QUAD__CH3_PIPE_TX_EQ_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RESET_BYP_HDSHK_CFG    32'h00000262
`define GTYE5_QUAD__CH3_RESET_BYP_HDSHK_CFG_SZ 32

`define GTYE5_QUAD__CH3_RESET_CFG    32'h00000263
`define GTYE5_QUAD__CH3_RESET_CFG_SZ 32

`define GTYE5_QUAD__CH3_RESET_LOOPER_ID_CFG    32'h00000264
`define GTYE5_QUAD__CH3_RESET_LOOPER_ID_CFG_SZ 32

`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG0    32'h00000265
`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG1    32'h00000266
`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG2    32'h00000267
`define GTYE5_QUAD__CH3_RESET_LOOP_ID_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RESET_TIME_CFG0    32'h00000268
`define GTYE5_QUAD__CH3_RESET_TIME_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RESET_TIME_CFG1    32'h00000269
`define GTYE5_QUAD__CH3_RESET_TIME_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RESET_TIME_CFG2    32'h0000026a
`define GTYE5_QUAD__CH3_RESET_TIME_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RESET_TIME_CFG3    32'h0000026b
`define GTYE5_QUAD__CH3_RESET_TIME_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RXOUTCLK_FREQ    32'h0000026c
`define GTYE5_QUAD__CH3_RXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH3_RXOUTCLK_REF_FREQ    32'h0000026d
`define GTYE5_QUAD__CH3_RXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH3_RXOUTCLK_REF_SOURCE    32'h0000026e
`define GTYE5_QUAD__CH3_RXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH3_RX_CDR_CFG0    32'h0000026f
`define GTYE5_QUAD__CH3_RX_CDR_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_CDR_CFG1    32'h00000270
`define GTYE5_QUAD__CH3_RX_CDR_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_CDR_CFG2    32'h00000271
`define GTYE5_QUAD__CH3_RX_CDR_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RX_CDR_CFG3    32'h00000272
`define GTYE5_QUAD__CH3_RX_CDR_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RX_CDR_CFG4    32'h00000273
`define GTYE5_QUAD__CH3_RX_CDR_CFG4_SZ 32

`define GTYE5_QUAD__CH3_RX_CRC_CFG0    32'h00000274
`define GTYE5_QUAD__CH3_RX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_CRC_CFG1    32'h00000275
`define GTYE5_QUAD__CH3_RX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_CRC_CFG2    32'h00000276
`define GTYE5_QUAD__CH3_RX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RX_CRC_CFG3    32'h00000277
`define GTYE5_QUAD__CH3_RX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RX_CTLE_CFG0    32'h00000278
`define GTYE5_QUAD__CH3_RX_CTLE_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_CTLE_CFG1    32'h00000279
`define GTYE5_QUAD__CH3_RX_CTLE_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_DACI2V_CFG0    32'h0000027a
`define GTYE5_QUAD__CH3_RX_DACI2V_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_DATA_RATE    32'h0000027b
`define GTYE5_QUAD__CH3_RX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH3_RX_DFE_CFG0    32'h0000027c
`define GTYE5_QUAD__CH3_RX_DFE_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG0    32'h0000027d
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG1    32'h0000027e
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG2    32'h0000027f
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG3    32'h00000280
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG4    32'h00000281
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG4_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG5    32'h00000282
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG5_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG6    32'h00000283
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG6_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG7    32'h00000284
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG7_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG8    32'h00000285
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG8_SZ 32

`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG9    32'h00000286
`define GTYE5_QUAD__CH3_RX_ELASTIC_BUF_CFG9_SZ 32

`define GTYE5_QUAD__CH3_RX_MISC_CFG0    32'h00000287
`define GTYE5_QUAD__CH3_RX_MISC_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_OOB_CFG0    32'h00000288
`define GTYE5_QUAD__CH3_RX_OOB_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_OOB_CFG1    32'h00000289
`define GTYE5_QUAD__CH3_RX_OOB_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_PAD_CFG0    32'h0000028a
`define GTYE5_QUAD__CH3_RX_PAD_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_PAD_CFG1    32'h0000028b
`define GTYE5_QUAD__CH3_RX_PAD_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_PCS_CFG0    32'h0000028c
`define GTYE5_QUAD__CH3_RX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_PCS_CFG1    32'h0000028d
`define GTYE5_QUAD__CH3_RX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_PCS_CFG2    32'h0000028e
`define GTYE5_QUAD__CH3_RX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RX_PCS_CFG3    32'h0000028f
`define GTYE5_QUAD__CH3_RX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RX_PCS_CFG4    32'h00000290
`define GTYE5_QUAD__CH3_RX_PCS_CFG4_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG0    32'h00000291
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG1    32'h00000292
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG2    32'h00000293
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG3    32'h00000294
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG4    32'h00000295
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG5    32'h00000296
`define GTYE5_QUAD__CH3_RX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH3_SIM_MODE    32'h00000297
`define GTYE5_QUAD__CH3_SIM_MODE_SZ 48

`define GTYE5_QUAD__CH3_SIM_RECEIVER_DETECT_PASS    32'h00000298
`define GTYE5_QUAD__CH3_SIM_RECEIVER_DETECT_PASS_SZ 40

`define GTYE5_QUAD__CH3_SIM_RESET_SPEEDUP    32'h00000299
`define GTYE5_QUAD__CH3_SIM_RESET_SPEEDUP_SZ 40

`define GTYE5_QUAD__CH3_SIM_TX_EIDLE_DRIVE_LEVEL    32'h0000029a
`define GTYE5_QUAD__CH3_SIM_TX_EIDLE_DRIVE_LEVEL_SZ 32

`define GTYE5_QUAD__CH3_TXOUTCLK_FREQ    32'h0000029b
`define GTYE5_QUAD__CH3_TXOUTCLK_FREQ_SZ 64

`define GTYE5_QUAD__CH3_TXOUTCLK_REF_FREQ    32'h0000029c
`define GTYE5_QUAD__CH3_TXOUTCLK_REF_FREQ_SZ 64

`define GTYE5_QUAD__CH3_TXOUTCLK_REF_SOURCE    32'h0000029d
`define GTYE5_QUAD__CH3_TXOUTCLK_REF_SOURCE_SZ 192

`define GTYE5_QUAD__CH3_TX_10G_CFG0    32'h0000029e
`define GTYE5_QUAD__CH3_TX_10G_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_10G_CFG1    32'h0000029f
`define GTYE5_QUAD__CH3_TX_10G_CFG1_SZ 32

`define GTYE5_QUAD__CH3_TX_10G_CFG2    32'h000002a0
`define GTYE5_QUAD__CH3_TX_10G_CFG2_SZ 32

`define GTYE5_QUAD__CH3_TX_10G_CFG3    32'h000002a1
`define GTYE5_QUAD__CH3_TX_10G_CFG3_SZ 32

`define GTYE5_QUAD__CH3_TX_ANA_CFG0    32'h000002a2
`define GTYE5_QUAD__CH3_TX_ANA_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_CRC_CFG0    32'h000002a3
`define GTYE5_QUAD__CH3_TX_CRC_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_CRC_CFG1    32'h000002a4
`define GTYE5_QUAD__CH3_TX_CRC_CFG1_SZ 32

`define GTYE5_QUAD__CH3_TX_CRC_CFG2    32'h000002a5
`define GTYE5_QUAD__CH3_TX_CRC_CFG2_SZ 32

`define GTYE5_QUAD__CH3_TX_CRC_CFG3    32'h000002a6
`define GTYE5_QUAD__CH3_TX_CRC_CFG3_SZ 32

`define GTYE5_QUAD__CH3_TX_DATA_RATE    32'h000002a7
`define GTYE5_QUAD__CH3_TX_DATA_RATE_SZ 64

`define GTYE5_QUAD__CH3_TX_DRV_CFG0    32'h000002a8
`define GTYE5_QUAD__CH3_TX_DRV_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_DRV_CFG1    32'h000002a9
`define GTYE5_QUAD__CH3_TX_DRV_CFG1_SZ 32

`define GTYE5_QUAD__CH3_TX_PCS_CFG0    32'h000002aa
`define GTYE5_QUAD__CH3_TX_PCS_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_PCS_CFG1    32'h000002ab
`define GTYE5_QUAD__CH3_TX_PCS_CFG1_SZ 32

`define GTYE5_QUAD__CH3_TX_PCS_CFG2    32'h000002ac
`define GTYE5_QUAD__CH3_TX_PCS_CFG2_SZ 32

`define GTYE5_QUAD__CH3_TX_PCS_CFG3    32'h000002ad
`define GTYE5_QUAD__CH3_TX_PCS_CFG3_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG0    32'h000002ae
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG0_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG1    32'h000002af
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG1_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG2    32'h000002b0
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG2_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG3    32'h000002b1
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG3_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG4    32'h000002b2
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG4_SZ 32

`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG5    32'h000002b3
`define GTYE5_QUAD__CH3_TX_PHALIGN_CFG5_SZ 32

`define GTYE5_QUAD__CH3_TX_PIPPM_CFG    32'h000002b4
`define GTYE5_QUAD__CH3_TX_PIPPM_CFG_SZ 32

`define GTYE5_QUAD__CH3_TX_SER_CFG0    32'h000002b5
`define GTYE5_QUAD__CH3_TX_SER_CFG0_SZ 32

`define GTYE5_QUAD__CHANNEL_CONNECTIVITY    32'h000002b6
`define GTYE5_QUAD__CHANNEL_CONNECTIVITY_SZ 32

`define GTYE5_QUAD__CTRL_RSV_CFG0    32'h000002b7
`define GTYE5_QUAD__CTRL_RSV_CFG0_SZ 32

`define GTYE5_QUAD__CTRL_RSV_CFG1    32'h000002b8
`define GTYE5_QUAD__CTRL_RSV_CFG1_SZ 32

`define GTYE5_QUAD__HS0_LCPLL_IPS_PIN_EN    32'h000002b9
`define GTYE5_QUAD__HS0_LCPLL_IPS_PIN_EN_SZ 1

`define GTYE5_QUAD__HS0_LCPLL_IPS_REFCLK_SEL    32'h000002ba
`define GTYE5_QUAD__HS0_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP0    32'h000002bb
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP0_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP1    32'h000002bc
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP1_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP2    32'h000002bd
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP2_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP3    32'h000002be
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP3_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP4    32'h000002bf
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP4_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP5    32'h000002c0
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP5_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP6    32'h000002c1
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP6_SZ 3

`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP7    32'h000002c2
`define GTYE5_QUAD__HS0_LCPLL_REFCLK_MAP7_SZ 3

`define GTYE5_QUAD__HS0_RPLL_IPS_PIN_EN    32'h000002c3
`define GTYE5_QUAD__HS0_RPLL_IPS_PIN_EN_SZ 1

`define GTYE5_QUAD__HS0_RPLL_IPS_REFCLK_SEL    32'h000002c4
`define GTYE5_QUAD__HS0_RPLL_IPS_REFCLK_SEL_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP0    32'h000002c5
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP0_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP1    32'h000002c6
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP1_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP2    32'h000002c7
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP2_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP3    32'h000002c8
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP3_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP4    32'h000002c9
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP4_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP5    32'h000002ca
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP5_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP6    32'h000002cb
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP6_SZ 3

`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP7    32'h000002cc
`define GTYE5_QUAD__HS0_RPLL_REFCLK_MAP7_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_IPS_PIN_EN    32'h000002cd
`define GTYE5_QUAD__HS1_LCPLL_IPS_PIN_EN_SZ 1

`define GTYE5_QUAD__HS1_LCPLL_IPS_REFCLK_SEL    32'h000002ce
`define GTYE5_QUAD__HS1_LCPLL_IPS_REFCLK_SEL_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP0    32'h000002cf
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP0_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP1    32'h000002d0
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP1_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP2    32'h000002d1
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP2_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP3    32'h000002d2
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP3_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP4    32'h000002d3
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP4_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP5    32'h000002d4
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP5_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP6    32'h000002d5
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP6_SZ 3

`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP7    32'h000002d6
`define GTYE5_QUAD__HS1_LCPLL_REFCLK_MAP7_SZ 3

`define GTYE5_QUAD__HS1_RPLL_IPS_PIN_EN    32'h000002d7
`define GTYE5_QUAD__HS1_RPLL_IPS_PIN_EN_SZ 1

`define GTYE5_QUAD__HS1_RPLL_IPS_REFCLK_SEL    32'h000002d8
`define GTYE5_QUAD__HS1_RPLL_IPS_REFCLK_SEL_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP0    32'h000002d9
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP0_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP1    32'h000002da
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP1_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP2    32'h000002db
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP2_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP3    32'h000002dc
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP3_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP4    32'h000002dd
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP4_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP5    32'h000002de
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP5_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP6    32'h000002df
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP6_SZ 3

`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP7    32'h000002e0
`define GTYE5_QUAD__HS1_RPLL_REFCLK_MAP7_SZ 3

`define GTYE5_QUAD__HSCLK0_HSDIST_CFG    32'h000002e1
`define GTYE5_QUAD__HSCLK0_HSDIST_CFG_SZ 32

`define GTYE5_QUAD__HSCLK0_INSTANTIATED    32'h000002e2
`define GTYE5_QUAD__HSCLK0_INSTANTIATED_SZ 1

`define GTYE5_QUAD__HSCLK0_LCPLL_CFG0    32'h000002e3
`define GTYE5_QUAD__HSCLK0_LCPLL_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK0_LCPLL_CFG1    32'h000002e4
`define GTYE5_QUAD__HSCLK0_LCPLL_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK0_LCPLL_CFG2    32'h000002e5
`define GTYE5_QUAD__HSCLK0_LCPLL_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG0    32'h000002e6
`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG1    32'h000002e7
`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG2    32'h000002e8
`define GTYE5_QUAD__HSCLK0_LCPLL_LGC_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_CFG0    32'h000002e9
`define GTYE5_QUAD__HSCLK0_RPLL_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_CFG1    32'h000002ea
`define GTYE5_QUAD__HSCLK0_RPLL_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_CFG2    32'h000002eb
`define GTYE5_QUAD__HSCLK0_RPLL_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG0    32'h000002ec
`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG1    32'h000002ed
`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG2    32'h000002ee
`define GTYE5_QUAD__HSCLK0_RPLL_LGC_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK0_RXRECCLK_SEL    32'h000002ef
`define GTYE5_QUAD__HSCLK0_RXRECCLK_SEL_SZ 2

`define GTYE5_QUAD__HSCLK1_HSDIST_CFG    32'h000002f0
`define GTYE5_QUAD__HSCLK1_HSDIST_CFG_SZ 32

`define GTYE5_QUAD__HSCLK1_INSTANTIATED    32'h000002f1
`define GTYE5_QUAD__HSCLK1_INSTANTIATED_SZ 1

`define GTYE5_QUAD__HSCLK1_LCPLL_CFG0    32'h000002f2
`define GTYE5_QUAD__HSCLK1_LCPLL_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK1_LCPLL_CFG1    32'h000002f3
`define GTYE5_QUAD__HSCLK1_LCPLL_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK1_LCPLL_CFG2    32'h000002f4
`define GTYE5_QUAD__HSCLK1_LCPLL_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG0    32'h000002f5
`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG1    32'h000002f6
`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG2    32'h000002f7
`define GTYE5_QUAD__HSCLK1_LCPLL_LGC_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_CFG0    32'h000002f8
`define GTYE5_QUAD__HSCLK1_RPLL_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_CFG1    32'h000002f9
`define GTYE5_QUAD__HSCLK1_RPLL_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_CFG2    32'h000002fa
`define GTYE5_QUAD__HSCLK1_RPLL_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG0    32'h000002fb
`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG0_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG1    32'h000002fc
`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG1_SZ 32

`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG2    32'h000002fd
`define GTYE5_QUAD__HSCLK1_RPLL_LGC_CFG2_SZ 32

`define GTYE5_QUAD__HSCLK1_RXRECCLK_SEL    32'h000002fe
`define GTYE5_QUAD__HSCLK1_RXRECCLK_SEL_SZ 2

`define GTYE5_QUAD__MEMORY_INIT_FILE    32'h000002ff
`define GTYE5_QUAD__MEMORY_INIT_FILE_SZ 32

`define GTYE5_QUAD__MST_RESET_CFG    32'h00000300
`define GTYE5_QUAD__MST_RESET_CFG_SZ 32

`define GTYE5_QUAD__PIN_CFG0    32'h00000301
`define GTYE5_QUAD__PIN_CFG0_SZ 32

`define GTYE5_QUAD__POR_CFG    32'h00000302
`define GTYE5_QUAD__POR_CFG_SZ 32

`define GTYE5_QUAD__QUAD_INSTANTIATED    32'h00000303
`define GTYE5_QUAD__QUAD_INSTANTIATED_SZ 1

`define GTYE5_QUAD__QUAD_SIM_MODE    32'h00000304
`define GTYE5_QUAD__QUAD_SIM_MODE_SZ 48

`define GTYE5_QUAD__QUAD_SIM_RESET_SPEEDUP    32'h00000305
`define GTYE5_QUAD__QUAD_SIM_RESET_SPEEDUP_SZ 40

`define GTYE5_QUAD__RCALBG0_CFG0    32'h00000306
`define GTYE5_QUAD__RCALBG0_CFG0_SZ 32

`define GTYE5_QUAD__RCALBG0_CFG1    32'h00000307
`define GTYE5_QUAD__RCALBG0_CFG1_SZ 32

`define GTYE5_QUAD__RCALBG0_CFG2    32'h00000308
`define GTYE5_QUAD__RCALBG0_CFG2_SZ 32

`define GTYE5_QUAD__RCALBG0_CFG3    32'h00000309
`define GTYE5_QUAD__RCALBG0_CFG3_SZ 32

`define GTYE5_QUAD__RCALBG0_CFG4    32'h0000030a
`define GTYE5_QUAD__RCALBG0_CFG4_SZ 32

`define GTYE5_QUAD__RCALBG0_CFG5    32'h0000030b
`define GTYE5_QUAD__RCALBG0_CFG5_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG0    32'h0000030c
`define GTYE5_QUAD__RCALBG1_CFG0_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG1    32'h0000030d
`define GTYE5_QUAD__RCALBG1_CFG1_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG2    32'h0000030e
`define GTYE5_QUAD__RCALBG1_CFG2_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG3    32'h0000030f
`define GTYE5_QUAD__RCALBG1_CFG3_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG4    32'h00000310
`define GTYE5_QUAD__RCALBG1_CFG4_SZ 32

`define GTYE5_QUAD__RCALBG1_CFG5    32'h00000311
`define GTYE5_QUAD__RCALBG1_CFG5_SZ 32

`define GTYE5_QUAD__RXRSTDONE_DIST_SEL    32'h00000312
`define GTYE5_QUAD__RXRSTDONE_DIST_SEL_SZ 32

`define GTYE5_QUAD__SIM_VERSION    32'h00000313
`define GTYE5_QUAD__SIM_VERSION_SZ 8

`define GTYE5_QUAD__STAT_NPI_REG_LIST    32'h00000314
`define GTYE5_QUAD__STAT_NPI_REG_LIST_SZ 32

`define GTYE5_QUAD__TERMPROG_CFG    32'h00000315
`define GTYE5_QUAD__TERMPROG_CFG_SZ 32

`define GTYE5_QUAD__TXRSTDONE_DIST_SEL    32'h00000316
`define GTYE5_QUAD__TXRSTDONE_DIST_SEL_SZ 32

`define GTYE5_QUAD__UB_CFG0    32'h00000317
`define GTYE5_QUAD__UB_CFG0_SZ 32

`endif  // B_GTYE5_QUAD_DEFINES_VH